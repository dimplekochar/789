-- VHDL global package produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
package ahir_system_global_package is -- 
  constant PJ_base_address : std_logic_vector(0 downto 0) := "0";
  constant ZJ_base_address : std_logic_vector(0 downto 0) := "0";
  constant a_base_address : std_logic_vector(3 downto 0) := "0000";
  constant image_base_address : std_logic_vector(3 downto 0) := "0000";
  constant kernel_base_address : std_logic_vector(3 downto 0) := "0000";
  constant mem_array_base_address : std_logic_vector(10 downto 0) := "00000000000";
  constant one_base_address : std_logic_vector(0 downto 0) := "0";
  constant total_base_address : std_logic_vector(0 downto 0) := "0";
  constant zer_base_address : std_logic_vector(0 downto 0) := "0";
  -- 
end package ahir_system_global_package;
