-- VHDL global package produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
package ahir_system_global_package is -- 
  constant mem_base_address : std_logic_vector(7 downto 0) := "00000000";
  constant next_pc1_base_address : std_logic_vector(0 downto 0) := "0";
  constant reg_base_address : std_logic_vector(7 downto 0) := "00000000";
  constant right_shift_base_address : std_logic_vector(0 downto 0) := "0";
  -- 
end package ahir_system_global_package;
