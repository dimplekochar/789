-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity accMemAccessDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    acc_mem_request : in  std_logic_vector(31 downto 0);
    acc_mem_responsel : out  std_logic_vector(31 downto 0);
    acc_mem_responseh : out  std_logic_vector(31 downto 0);
    accessMem_call_reqs : out  std_logic_vector(0 downto 0);
    accessMem_call_acks : in   std_logic_vector(0 downto 0);
    accessMem_call_data : out  std_logic_vector(28 downto 0);
    accessMem_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMem_return_reqs : out  std_logic_vector(0 downto 0);
    accessMem_return_acks : in   std_logic_vector(0 downto 0);
    accessMem_return_data : in   std_logic_vector(63 downto 0);
    accessMem_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accMemAccessDaemon;
architecture accMemAccessDaemon_arch of accMemAccessDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal acc_mem_request_buffer :  std_logic_vector(31 downto 0);
  signal acc_mem_request_update_enable: Boolean;
  -- output port buffer signals
  signal acc_mem_responsel_buffer :  std_logic_vector(31 downto 0);
  signal acc_mem_responsel_update_enable: Boolean;
  signal acc_mem_responseh_buffer :  std_logic_vector(31 downto 0);
  signal acc_mem_responseh_update_enable: Boolean;
  signal accMemAccessDaemon_CP_491_start: Boolean;
  signal accMemAccessDaemon_CP_491_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(11 downto 0);
      write_data : in  std_logic_vector(15 downto 0);
      read_datal : out  std_logic_vector(63 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_127_call_ack_1 : boolean;
  signal call_stmt_127_call_req_1 : boolean;
  signal W_acc_mem_responsel_136_inst_ack_1 : boolean;
  signal W_acc_mem_responsel_136_inst_req_1 : boolean;
  signal W_acc_mem_responsel_136_inst_ack_0 : boolean;
  signal W_acc_mem_responseh_139_inst_ack_1 : boolean;
  signal W_acc_mem_responseh_139_inst_ack_0 : boolean;
  signal W_acc_mem_responsel_136_inst_req_0 : boolean;
  signal W_acc_mem_responseh_139_inst_req_1 : boolean;
  signal W_acc_mem_responseh_139_inst_req_0 : boolean;
  signal W_cmd_108_inst_req_0 : boolean;
  signal W_cmd_108_inst_ack_0 : boolean;
  signal W_cmd_108_inst_req_1 : boolean;
  signal W_cmd_108_inst_ack_1 : boolean;
  signal call_stmt_127_call_req_0 : boolean;
  signal call_stmt_127_call_ack_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accMemAccessDaemon_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 32) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= acc_mem_request;
  acc_mem_request_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(tag_length + 31 downto 32) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 31 downto 32);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accMemAccessDaemon_CP_491_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accMemAccessDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= acc_mem_responsel_buffer;
  acc_mem_responsel <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(63 downto 32) <= acc_mem_responseh_buffer;
  acc_mem_responseh <= out_buffer_data_out(63 downto 32);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accMemAccessDaemon_CP_491_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accMemAccessDaemon_CP_491_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accMemAccessDaemon_CP_491_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,accMemAccessDaemon_CP_491_start,"accMemAccessDaemon cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,accMemAccessDaemon_CP_491_symbol, "accMemAccessDaemon cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accMemAccessDaemon_CP_491: Block -- control-path 
    signal accMemAccessDaemon_CP_491_elements: BooleanArray(9 downto 0);
    -- 
  begin -- 
    accMemAccessDaemon_CP_491_elements(0) <= accMemAccessDaemon_CP_491_start;
    accMemAccessDaemon_CP_491_symbol <= accMemAccessDaemon_CP_491_elements(9);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (17) 
      -- CP-element group 0: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_141_update_start_
      -- CP-element group 0: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_138_update_start_
      -- CP-element group 0: 	 assign_stmt_110_to_assign_stmt_141/call_stmt_127_Update/ccr
      -- CP-element group 0: 	 assign_stmt_110_to_assign_stmt_141/call_stmt_127_Update/$entry
      -- CP-element group 0: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_138_Update/req
      -- CP-element group 0: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_138_Update/$entry
      -- CP-element group 0: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_141_Update/$entry
      -- CP-element group 0: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_141_Update/req
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_110_to_assign_stmt_141/$entry
      -- CP-element group 0: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_110_sample_start_
      -- CP-element group 0: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_110_update_start_
      -- CP-element group 0: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_110_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_110_Sample/req
      -- CP-element group 0: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_110_Update/$entry
      -- CP-element group 0: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_110_Update/req
      -- CP-element group 0: 	 assign_stmt_110_to_assign_stmt_141/call_stmt_127_update_start_
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_491_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_491_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_491_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:W_cmd_108_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:W_cmd_108_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:W_acc_mem_responseh_139_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:call_stmt_127_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:W_acc_mem_responsel_136_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accMemAccessDaemon_CP_491_elements(0), ack => W_cmd_108_inst_req_0); -- 
    req_509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accMemAccessDaemon_CP_491_elements(0), ack => W_cmd_108_inst_req_1); -- 
    req_551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accMemAccessDaemon_CP_491_elements(0), ack => W_acc_mem_responseh_139_inst_req_1); -- 
    ccr_523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accMemAccessDaemon_CP_491_elements(0), ack => call_stmt_127_call_req_1); -- 
    req_537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accMemAccessDaemon_CP_491_elements(0), ack => W_acc_mem_responsel_136_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_110_sample_completed_
      -- CP-element group 1: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_110_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_110_Sample/ack
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_491_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_491_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_491_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:W_cmd_108_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_cmd_108_inst_ack_0, ack => accMemAccessDaemon_CP_491_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_110_update_completed_
      -- CP-element group 2: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_110_Update/$exit
      -- CP-element group 2: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_110_Update/ack
      -- CP-element group 2: 	 assign_stmt_110_to_assign_stmt_141/call_stmt_127_sample_start_
      -- CP-element group 2: 	 assign_stmt_110_to_assign_stmt_141/call_stmt_127_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_110_to_assign_stmt_141/call_stmt_127_Sample/crr
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_491_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_491_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_491_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:W_cmd_108_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:call_stmt_127_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_cmd_108_inst_ack_1, ack => accMemAccessDaemon_CP_491_elements(2)); -- 
    crr_518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accMemAccessDaemon_CP_491_elements(2), ack => call_stmt_127_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_110_to_assign_stmt_141/call_stmt_127_sample_completed_
      -- CP-element group 3: 	 assign_stmt_110_to_assign_stmt_141/call_stmt_127_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_110_to_assign_stmt_141/call_stmt_127_Sample/cra
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_491_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_491_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_491_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:call_stmt_127_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_127_call_ack_0, ack => accMemAccessDaemon_CP_491_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_138_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_138_sample_start_
      -- CP-element group 4: 	 assign_stmt_110_to_assign_stmt_141/call_stmt_127_Update/cca
      -- CP-element group 4: 	 assign_stmt_110_to_assign_stmt_141/call_stmt_127_Update/$exit
      -- CP-element group 4: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_141_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_141_sample_start_
      -- CP-element group 4: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_138_Sample/req
      -- CP-element group 4: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_141_Sample/req
      -- CP-element group 4: 	 assign_stmt_110_to_assign_stmt_141/call_stmt_127_update_completed_
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_491_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_491_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_491_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:call_stmt_127_call_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:W_acc_mem_responseh_139_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:W_acc_mem_responsel_136_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    cca_524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_127_call_ack_1, ack => accMemAccessDaemon_CP_491_elements(4)); -- 
    req_546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accMemAccessDaemon_CP_491_elements(4), ack => W_acc_mem_responseh_139_inst_req_0); -- 
    req_532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accMemAccessDaemon_CP_491_elements(4), ack => W_acc_mem_responsel_136_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_138_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_138_sample_completed_
      -- CP-element group 5: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_138_Sample/ack
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_491_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_491_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_491_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:W_acc_mem_responsel_136_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc_mem_responsel_136_inst_ack_0, ack => accMemAccessDaemon_CP_491_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_138_Update/$exit
      -- CP-element group 6: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_138_update_completed_
      -- CP-element group 6: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_138_Update/ack
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_491_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_491_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_491_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:W_acc_mem_responsel_136_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc_mem_responsel_136_inst_ack_1, ack => accMemAccessDaemon_CP_491_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_141_Sample/$exit
      -- CP-element group 7: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_141_sample_completed_
      -- CP-element group 7: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_141_Sample/ack
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_491_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_491_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_491_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:W_acc_mem_responseh_139_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc_mem_responseh_139_inst_ack_0, ack => accMemAccessDaemon_CP_491_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_141_update_completed_
      -- CP-element group 8: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_141_Update/$exit
      -- CP-element group 8: 	 assign_stmt_110_to_assign_stmt_141/assign_stmt_141_Update/ack
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_491_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_491_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_491_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:W_acc_mem_responseh_139_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc_mem_responseh_139_inst_ack_1, ack => accMemAccessDaemon_CP_491_elements(8)); -- 
    -- CP-element group 9:  join  transition  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 $exit
      -- CP-element group 9: 	 assign_stmt_110_to_assign_stmt_141/$exit
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_491_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_491_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_491_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    accMemAccessDaemon_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "accMemAccessDaemon_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accMemAccessDaemon_CP_491_elements(6) & accMemAccessDaemon_CP_491_elements(8);
      gj_accMemAccessDaemon_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accMemAccessDaemon_CP_491_elements(9), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal addr_122 : std_logic_vector(11 downto 0);
    signal cmd_110 : std_logic_vector(31 downto 0);
    signal rdata0_135 : std_logic_vector(31 downto 0);
    signal rdata1_131 : std_logic_vector(31 downto 0);
    signal rdatal_127 : std_logic_vector(63 downto 0);
    signal rwbar_114 : std_logic_vector(0 downto 0);
    signal wdata_118 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    -- logger for split-operator slice_113_inst flow-through 
    process(rwbar_114) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:slice_113_inst:flowthrough inputs: " & " cmd_110 = "& Convert_SLV_To_Hex_String(cmd_110) & " outputs:" & " rwbar_114= "  & Convert_SLV_To_Hex_String(rwbar_114));
      --
    end process; 
    -- flow-through slice operator slice_113_inst
    rwbar_114 <= cmd_110(31 downto 31);
    -- logger for split-operator slice_117_inst flow-through 
    process(wdata_118) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:slice_117_inst:flowthrough inputs: " & " cmd_110 = "& Convert_SLV_To_Hex_String(cmd_110) & " outputs:" & " wdata_118= "  & Convert_SLV_To_Hex_String(wdata_118));
      --
    end process; 
    -- flow-through slice operator slice_117_inst
    wdata_118 <= cmd_110(27 downto 12);
    -- logger for split-operator slice_121_inst flow-through 
    process(addr_122) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:slice_121_inst:flowthrough inputs: " & " cmd_110 = "& Convert_SLV_To_Hex_String(cmd_110) & " outputs:" & " addr_122= "  & Convert_SLV_To_Hex_String(addr_122));
      --
    end process; 
    -- flow-through slice operator slice_121_inst
    addr_122 <= cmd_110(11 downto 0);
    -- logger for split-operator slice_130_inst flow-through 
    process(rdata1_131) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:slice_130_inst:flowthrough inputs: " & " rdatal_127 = "& Convert_SLV_To_Hex_String(rdatal_127) & " outputs:" & " rdata1_131= "  & Convert_SLV_To_Hex_String(rdata1_131));
      --
    end process; 
    -- flow-through slice operator slice_130_inst
    rdata1_131 <= rdatal_127(63 downto 32);
    -- logger for split-operator slice_134_inst flow-through 
    process(rdata0_135) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:slice_134_inst:flowthrough inputs: " & " rdatal_127 = "& Convert_SLV_To_Hex_String(rdatal_127) & " outputs:" & " rdata0_135= "  & Convert_SLV_To_Hex_String(rdata0_135));
      --
    end process; 
    -- flow-through slice operator slice_134_inst
    rdata0_135 <= rdatal_127(31 downto 0);
    -- logger for split-operator W_acc_mem_responseh_139_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_acc_mem_responseh_139_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:W_acc_mem_responseh_139_inst:started:   inputs: " & " rdata1_131 = "& Convert_SLV_To_Hex_String(rdata1_131));
          --
        end if; 
        if W_acc_mem_responseh_139_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:W_acc_mem_responseh_139_inst:finished:  outputs: " & " acc_mem_responseh_buffer= "  & Convert_SLV_To_Hex_String(acc_mem_responseh_buffer));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_acc_mem_responseh_139_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_acc_mem_responseh_139_inst_req_0;
      W_acc_mem_responseh_139_inst_ack_0<= wack(0);
      rreq(0) <= W_acc_mem_responseh_139_inst_req_1;
      W_acc_mem_responseh_139_inst_ack_1<= rack(0);
      W_acc_mem_responseh_139_inst : InterlockBuffer generic map ( -- 
        name => "W_acc_mem_responseh_139_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rdata1_131,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => acc_mem_responseh_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_acc_mem_responsel_136_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_acc_mem_responsel_136_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:W_acc_mem_responsel_136_inst:started:   inputs: " & " rdata0_135 = "& Convert_SLV_To_Hex_String(rdata0_135));
          --
        end if; 
        if W_acc_mem_responsel_136_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:W_acc_mem_responsel_136_inst:finished:  outputs: " & " acc_mem_responsel_buffer= "  & Convert_SLV_To_Hex_String(acc_mem_responsel_buffer));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_acc_mem_responsel_136_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_acc_mem_responsel_136_inst_req_0;
      W_acc_mem_responsel_136_inst_ack_0<= wack(0);
      rreq(0) <= W_acc_mem_responsel_136_inst_req_1;
      W_acc_mem_responsel_136_inst_ack_1<= rack(0);
      W_acc_mem_responsel_136_inst : InterlockBuffer generic map ( -- 
        name => "W_acc_mem_responsel_136_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rdata0_135,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => acc_mem_responsel_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_cmd_108_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_cmd_108_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:W_cmd_108_inst:started:   inputs: " & " acc_mem_request_buffer = "& Convert_SLV_To_Hex_String(acc_mem_request_buffer));
          --
        end if; 
        if W_cmd_108_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:W_cmd_108_inst:finished:  outputs: " & " cmd_110= "  & Convert_SLV_To_Hex_String(cmd_110));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_cmd_108_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_cmd_108_inst_req_0;
      W_cmd_108_inst_ack_0<= wack(0);
      rreq(0) <= W_cmd_108_inst_req_1;
      W_cmd_108_inst_ack_1<= rack(0);
      W_cmd_108_inst : InterlockBuffer generic map ( -- 
        name => "W_cmd_108_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_mem_request_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => cmd_110,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator call_stmt_127_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_127_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:call_stmt_127_call:started:  Call to module accessMem inputs: " & " rwbar_114 = "& Convert_SLV_To_Hex_String(rwbar_114) & " addr_122 = "& Convert_SLV_To_Hex_String(addr_122) & " wdata_118 = "& Convert_SLV_To_Hex_String(wdata_118));
          --
        end if; 
        if call_stmt_127_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:call_stmt_127_call:finished:  outputs: " & " rdatal_127= "  & Convert_SLV_To_Hex_String(rdatal_127));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_127_call 
    accessMem_call_group_0: Block -- 
      signal data_in: std_logic_vector(28 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_127_call_req_0;
      call_stmt_127_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_127_call_req_1;
      call_stmt_127_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMem_call_group_0_gI: SplitGuardInterface generic map(name => "accessMem_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rwbar_114 & addr_122 & wdata_118;
      rdatal_127 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 29,
        owidth => 29,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMem_call_reqs(0),
          ackR => accessMem_call_acks(0),
          dataR => accessMem_call_data(28 downto 0),
          tagR => accessMem_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMem_return_acks(0), -- cross-over
          ackL => accessMem_return_reqs(0), -- cross-over
          dataL => accessMem_return_data(63 downto 0),
          tagL => accessMem_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end accMemAccessDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity accessMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    read_write_bar : in  std_logic_vector(0 downto 0);
    addr : in  std_logic_vector(11 downto 0);
    write_data : in  std_logic_vector(15 downto 0);
    read_datal : out  std_logic_vector(63 downto 0);
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(10 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessMem;
architecture accessMem_arch of accessMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 29)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal read_write_bar_buffer :  std_logic_vector(0 downto 0);
  signal read_write_bar_update_enable: Boolean;
  signal addr_buffer :  std_logic_vector(11 downto 0);
  signal addr_update_enable: Boolean;
  signal write_data_buffer :  std_logic_vector(15 downto 0);
  signal write_data_update_enable: Boolean;
  -- output port buffer signals
  signal read_datal_buffer :  std_logic_vector(63 downto 0);
  signal read_datal_update_enable: Boolean;
  signal accessMem_CP_0_start: Boolean;
  signal accessMem_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_28_load_0_req_0 : boolean;
  signal array_obj_ref_28_load_0_ack_0 : boolean;
  signal array_obj_ref_28_load_0_req_1 : boolean;
  signal array_obj_ref_28_load_0_ack_1 : boolean;
  signal ADD_u12_u12_34_inst_req_0 : boolean;
  signal ADD_u12_u12_34_inst_ack_0 : boolean;
  signal ADD_u12_u12_34_inst_req_1 : boolean;
  signal ADD_u12_u12_34_inst_ack_1 : boolean;
  signal W_read_write_bar_36_delayed_1_0_36_inst_req_0 : boolean;
  signal W_read_write_bar_36_delayed_1_0_36_inst_ack_0 : boolean;
  signal W_read_write_bar_36_delayed_1_0_36_inst_req_1 : boolean;
  signal W_read_write_bar_36_delayed_1_0_36_inst_ack_1 : boolean;
  signal array_obj_ref_42_load_0_req_0 : boolean;
  signal array_obj_ref_42_load_0_ack_0 : boolean;
  signal array_obj_ref_42_load_0_req_1 : boolean;
  signal array_obj_ref_42_load_0_ack_1 : boolean;
  signal ADD_u12_u12_48_inst_req_0 : boolean;
  signal ADD_u12_u12_48_inst_ack_0 : boolean;
  signal ADD_u12_u12_48_inst_req_1 : boolean;
  signal ADD_u12_u12_48_inst_ack_1 : boolean;
  signal W_read_write_bar_47_delayed_1_0_50_inst_req_0 : boolean;
  signal W_read_write_bar_47_delayed_1_0_50_inst_ack_0 : boolean;
  signal W_read_write_bar_47_delayed_1_0_50_inst_req_1 : boolean;
  signal W_read_write_bar_47_delayed_1_0_50_inst_ack_1 : boolean;
  signal array_obj_ref_56_load_0_req_0 : boolean;
  signal array_obj_ref_56_load_0_ack_0 : boolean;
  signal array_obj_ref_56_load_0_req_1 : boolean;
  signal array_obj_ref_56_load_0_ack_1 : boolean;
  signal ADD_u12_u12_62_inst_req_0 : boolean;
  signal ADD_u12_u12_62_inst_ack_0 : boolean;
  signal ADD_u12_u12_62_inst_req_1 : boolean;
  signal ADD_u12_u12_62_inst_ack_1 : boolean;
  signal W_read_write_bar_58_delayed_1_0_64_inst_req_0 : boolean;
  signal W_read_write_bar_58_delayed_1_0_64_inst_ack_0 : boolean;
  signal W_read_write_bar_58_delayed_1_0_64_inst_req_1 : boolean;
  signal W_read_write_bar_58_delayed_1_0_64_inst_ack_1 : boolean;
  signal array_obj_ref_70_load_0_req_0 : boolean;
  signal array_obj_ref_70_load_0_ack_0 : boolean;
  signal array_obj_ref_70_load_0_req_1 : boolean;
  signal array_obj_ref_70_load_0_ack_1 : boolean;
  signal W_t_read_data0_69_delayed_1_0_72_inst_req_0 : boolean;
  signal W_t_read_data0_69_delayed_1_0_72_inst_ack_0 : boolean;
  signal W_t_read_data0_69_delayed_1_0_72_inst_req_1 : boolean;
  signal W_t_read_data0_69_delayed_1_0_72_inst_ack_1 : boolean;
  signal W_read_write_bar_63_delayed_6_0_75_inst_req_0 : boolean;
  signal W_read_write_bar_63_delayed_6_0_75_inst_ack_0 : boolean;
  signal W_read_write_bar_63_delayed_6_0_75_inst_req_1 : boolean;
  signal W_read_write_bar_63_delayed_6_0_75_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_86_inst_req_0 : boolean;
  signal CONCAT_u32_u64_86_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_86_inst_req_1 : boolean;
  signal CONCAT_u32_u64_86_inst_ack_1 : boolean;
  signal array_obj_ref_90_store_0_req_0 : boolean;
  signal array_obj_ref_90_store_0_ack_0 : boolean;
  signal array_obj_ref_90_store_0_req_1 : boolean;
  signal array_obj_ref_90_store_0_ack_1 : boolean;
  signal W_read_write_bar_79_delayed_7_0_93_inst_req_0 : boolean;
  signal W_read_write_bar_79_delayed_7_0_93_inst_ack_0 : boolean;
  signal W_read_write_bar_79_delayed_7_0_93_inst_req_1 : boolean;
  signal W_read_write_bar_79_delayed_7_0_93_inst_ack_1 : boolean;
  signal MUX_100_inst_req_0 : boolean;
  signal MUX_100_inst_ack_0 : boolean;
  signal MUX_100_inst_req_1 : boolean;
  signal MUX_100_inst_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessMem_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 29) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= read_write_bar;
  read_write_bar_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(12 downto 1) <= addr;
  addr_buffer <= in_buffer_data_out(12 downto 1);
  in_buffer_data_in(28 downto 13) <= write_data;
  write_data_buffer <= in_buffer_data_out(28 downto 13);
  in_buffer_data_in(tag_length + 28 downto 29) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 28 downto 29);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 4) := (0 => 14,1 => 14,2 => 14,3 => 1,4 => 14);
    constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 14);
    constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 5); -- 
  begin -- 
    preds <= read_write_bar_update_enable & addr_update_enable & write_data_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessMem_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= read_datal_buffer;
  read_datal <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 14,1 => 1,2 => 14);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMem_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  read_datal_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 29) := "read_datal_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_read_datal_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => read_datal_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 14,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 14,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessMem_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 14,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMem_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,accessMem_CP_0_start,"accessMem cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,accessMem_CP_0_symbol, "accessMem cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessMem_CP_0: Block -- control-path 
    signal accessMem_CP_0_elements: BooleanArray(79 downto 0);
    -- 
  begin -- 
    accessMem_CP_0_elements(0) <= accessMem_CP_0_start;
    accessMem_CP_0_symbol <= accessMem_CP_0_elements(79);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- logger for CP element group accessMem_CP_0_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	22 
    -- CP-element group 1: 	26 
    -- CP-element group 1: 	34 
    -- CP-element group 1: 	38 
    -- CP-element group 1: 	6 
    -- CP-element group 1: 	10 
    -- CP-element group 1: 	14 
    -- CP-element group 1: 	50 
    -- CP-element group 1: 	58 
    -- CP-element group 1: 	62 
    -- CP-element group 1:  members (53) 
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/$entry
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_word_address_calculated
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_root_address_calculated
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_offset_calculated
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_index_resized_0
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_index_scaled_0
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_index_computed_0
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_index_resize_0/$entry
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_index_resize_0/$exit
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_index_resize_0/index_resize_req
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_index_resize_0/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_index_scale_0/$entry
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_index_scale_0/$exit
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_index_scale_0/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_index_scale_0/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_final_index_sum_regn/$entry
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_final_index_sum_regn/$exit
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_final_index_sum_regn/req
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_final_index_sum_regn/ack
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_base_plus_offset/$entry
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_base_plus_offset/$exit
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_base_plus_offset/sum_rename_req
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_base_plus_offset/sum_rename_ack
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_word_addrgen/$entry
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_word_addrgen/$exit
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_word_addrgen/root_register_req
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_word_addrgen/root_register_ack
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_word_address_calculated
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_root_address_calculated
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_offset_calculated
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_index_resized_0
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_index_scaled_0
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_index_computed_0
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_index_resize_0/$entry
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_index_resize_0/$exit
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_index_resize_0/index_resize_req
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_index_resize_0/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_index_scale_0/$entry
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_index_scale_0/$exit
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_index_scale_0/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_index_scale_0/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_final_index_sum_regn/$entry
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_final_index_sum_regn/$exit
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_final_index_sum_regn/req
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_final_index_sum_regn/ack
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_base_plus_offset/$entry
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_base_plus_offset/$exit
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_base_plus_offset/sum_rename_req
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_base_plus_offset/sum_rename_ack
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_word_addrgen/$entry
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_word_addrgen/$exit
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_word_addrgen/root_register_req
      -- CP-element group 1: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_CP_0_elements(1) <= accessMem_CP_0_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	36 
    -- CP-element group 2: 	40 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	52 
    -- CP-element group 2: 	60 
    -- CP-element group 2: 	64 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	75 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_29_to_assign_stmt_101/read_write_bar_update_enable
      -- CP-element group 2: 	 assign_stmt_29_to_assign_stmt_101/read_write_bar_update_enable_out
      -- 
    -- logger for CP element group accessMem_CP_0_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 28) := "accessMem_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(24) & accessMem_CP_0_elements(28) & accessMem_CP_0_elements(36) & accessMem_CP_0_elements(40) & accessMem_CP_0_elements(16) & accessMem_CP_0_elements(8) & accessMem_CP_0_elements(12) & accessMem_CP_0_elements(52) & accessMem_CP_0_elements(60) & accessMem_CP_0_elements(64);
      gj_accessMem_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	24 
    -- CP-element group 3: 	36 
    -- CP-element group 3: 	8 
    -- CP-element group 3: 	12 
    -- CP-element group 3: 	60 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	76 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_29_to_assign_stmt_101/addr_update_enable
      -- CP-element group 3: 	 assign_stmt_29_to_assign_stmt_101/addr_update_enable_out
      -- 
    -- logger for CP element group accessMem_CP_0_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "accessMem_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(24) & accessMem_CP_0_elements(36) & accessMem_CP_0_elements(8) & accessMem_CP_0_elements(12) & accessMem_CP_0_elements(60);
      gj_accessMem_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	60 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	77 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_29_to_assign_stmt_101/write_data_update_enable
      -- CP-element group 4: 	 assign_stmt_29_to_assign_stmt_101/write_data_update_enable_out
      -- 
    -- logger for CP element group accessMem_CP_0_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "accessMem_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMem_CP_0_elements(60);
      gj_accessMem_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	78 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	67 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_29_to_assign_stmt_101/read_datal_update_enable
      -- CP-element group 5: 	 assign_stmt_29_to_assign_stmt_101/read_datal_update_enable_in
      -- 
    -- logger for CP element group accessMem_CP_0_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_CP_0_elements(5) <= accessMem_CP_0_elements(78);
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	1 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	8 
    -- CP-element group 6: 	60 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (5) 
      -- CP-element group 6: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_sample_start_
      -- CP-element group 6: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_Sample/$entry
      -- CP-element group 6: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_Sample/word_access_start/$entry
      -- CP-element group 6: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_Sample/word_access_start/word_0/$entry
      -- CP-element group 6: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_28_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_59_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_59_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(6), ack => array_obj_ref_28_load_0_req_0); -- 
    accessMem_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 14,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 28) := "accessMem_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(8) & accessMem_CP_0_elements(60);
      gj_accessMem_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: marked-predecessors 
    -- CP-element group 7: 	9 
    -- CP-element group 7: 	48 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	9 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_update_start_
      -- CP-element group 7: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_Update/$entry
      -- CP-element group 7: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_Update/word_access_complete/$entry
      -- CP-element group 7: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_Update/word_access_complete/word_0/$entry
      -- CP-element group 7: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_28_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_70_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_70_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(7), ack => array_obj_ref_28_load_0_req_1); -- 
    accessMem_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "accessMem_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(9) & accessMem_CP_0_elements(48);
      gj_accessMem_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	70 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: 	3 
    -- CP-element group 8: 	6 
    -- CP-element group 8:  members (5) 
      -- CP-element group 8: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_sample_completed_
      -- CP-element group 8: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_Sample/$exit
      -- CP-element group 8: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_Sample/word_access_start/$exit
      -- CP-element group 8: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_Sample/word_access_start/word_0/$exit
      -- CP-element group 8: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group accessMem_CP_0_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_28_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_60_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_28_load_0_ack_0, ack => accessMem_CP_0_elements(8)); -- 
    -- CP-element group 9:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	7 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	46 
    -- CP-element group 9: marked-successors 
    -- CP-element group 9: 	7 
    -- CP-element group 9:  members (9) 
      -- CP-element group 9: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_update_completed_
      -- CP-element group 9: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_Update/$exit
      -- CP-element group 9: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_Update/word_access_complete/$exit
      -- CP-element group 9: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_Update/word_access_complete/word_0/$exit
      -- CP-element group 9: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_Update/word_access_complete/word_0/ca
      -- CP-element group 9: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_Update/array_obj_ref_28_Merge/$entry
      -- CP-element group 9: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_Update/array_obj_ref_28_Merge/$exit
      -- CP-element group 9: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_Update/array_obj_ref_28_Merge/merge_req
      -- CP-element group 9: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_Update/array_obj_ref_28_Merge/merge_ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(9) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_28_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_71_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_28_load_0_ack_1, ack => accessMem_CP_0_elements(9)); -- 
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	1 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_34_sample_start_
      -- CP-element group 10: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_34_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_34_Sample/rr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:ADD_u12_u12_34_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_84_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_84_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(10), ack => ADD_u12_u12_34_inst_req_0); -- 
    accessMem_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 14,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(12);
      gj_accessMem_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	20 
    -- CP-element group 11: 	13 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_34_update_start_
      -- CP-element group 11: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_34_Update/$entry
      -- CP-element group 11: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_34_Update/cr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:ADD_u12_u12_34_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_89_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_89_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(11), ack => ADD_u12_u12_34_inst_req_1); -- 
    accessMem_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(20) & accessMem_CP_0_elements(13);
      gj_accessMem_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: 	3 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_34_sample_completed_
      -- CP-element group 12: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_34_Sample/$exit
      -- CP-element group 12: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_34_Sample/ra
      -- 
    -- logger for CP element group accessMem_CP_0_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:ADD_u12_u12_34_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_85_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_34_inst_ack_0, ack => accessMem_CP_0_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	18 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	11 
    -- CP-element group 13:  members (29) 
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_offset_calculated
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_index_resized_0
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_index_scaled_0
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_index_computed_0
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_index_resize_0/$entry
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_index_resize_0/$exit
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_index_resize_0/index_resize_req
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_34_update_completed_
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_34_Update/$exit
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_34_Update/ca
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_word_address_calculated
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_root_address_calculated
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_index_resize_0/index_resize_ack
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_index_scale_0/$entry
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_index_scale_0/$exit
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_index_scale_0/scale_rename_req
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_index_scale_0/scale_rename_ack
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_final_index_sum_regn/$entry
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_final_index_sum_regn/$exit
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_final_index_sum_regn/req
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_final_index_sum_regn/ack
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_base_plus_offset/$entry
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_base_plus_offset/$exit
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_base_plus_offset/sum_rename_req
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_base_plus_offset/sum_rename_ack
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_word_addrgen/$entry
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_word_addrgen/$exit
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_word_addrgen/root_register_req
      -- CP-element group 13: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:ADD_u12_u12_34_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_90_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_34_inst_ack_1, ack => accessMem_CP_0_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	1 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_38_sample_start_
      -- CP-element group 14: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_38_Sample/$entry
      -- CP-element group 14: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_38_Sample/req
      -- 
    -- logger for CP element group accessMem_CP_0_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_36_delayed_1_0_36_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_98_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_98_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(14), ack => W_read_write_bar_36_delayed_1_0_36_inst_req_0); -- 
    accessMem_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 14,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(16);
      gj_accessMem_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	20 
    -- CP-element group 15: 	17 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_38_update_start_
      -- CP-element group 15: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_38_Update/$entry
      -- CP-element group 15: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_38_Update/req
      -- 
    -- logger for CP element group accessMem_CP_0_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_36_delayed_1_0_36_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(15), ack => W_read_write_bar_36_delayed_1_0_36_inst_req_1); -- 
    accessMem_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(20) & accessMem_CP_0_elements(17);
      gj_accessMem_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_38_sample_completed_
      -- CP-element group 16: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_38_Sample/$exit
      -- CP-element group 16: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_38_Sample/ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_36_delayed_1_0_36_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_99_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_36_delayed_1_0_36_inst_ack_0, ack => accessMem_CP_0_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	15 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_38_update_completed_
      -- CP-element group 17: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_38_Update/$exit
      -- CP-element group 17: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_38_Update/ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_36_delayed_1_0_36_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_36_delayed_1_0_36_inst_ack_1, ack => accessMem_CP_0_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: 	13 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: 	60 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (5) 
      -- CP-element group 18: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_sample_start_
      -- CP-element group 18: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_Sample/$entry
      -- CP-element group 18: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_Sample/word_access_start/$entry
      -- CP-element group 18: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_Sample/word_access_start/word_0/$entry
      -- CP-element group 18: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_42_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(18), ack => array_obj_ref_42_load_0_req_0); -- 
    accessMem_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(17) & accessMem_CP_0_elements(13) & accessMem_CP_0_elements(20) & accessMem_CP_0_elements(60);
      gj_accessMem_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	21 
    -- CP-element group 19: 	56 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_update_start_
      -- CP-element group 19: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_Update/$entry
      -- CP-element group 19: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_Update/word_access_complete/$entry
      -- CP-element group 19: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_Update/word_access_complete/word_0/$entry
      -- CP-element group 19: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_42_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(19), ack => array_obj_ref_42_load_0_req_1); -- 
    accessMem_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(21) & accessMem_CP_0_elements(56);
      gj_accessMem_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	71 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: 	11 
    -- CP-element group 20: 	15 
    -- CP-element group 20:  members (5) 
      -- CP-element group 20: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_sample_completed_
      -- CP-element group 20: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_Sample/$exit
      -- CP-element group 20: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_Sample/word_access_start/$exit
      -- CP-element group 20: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_Sample/word_access_start/word_0/$exit
      -- CP-element group 20: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group accessMem_CP_0_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_42_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_42_load_0_ack_0, ack => accessMem_CP_0_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	54 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	19 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_update_completed_
      -- CP-element group 21: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_Update/$exit
      -- CP-element group 21: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_Update/word_access_complete/$exit
      -- CP-element group 21: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_Update/word_access_complete/word_0/$exit
      -- CP-element group 21: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_Update/word_access_complete/word_0/ca
      -- CP-element group 21: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_Update/array_obj_ref_42_Merge/$entry
      -- CP-element group 21: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_Update/array_obj_ref_42_Merge/$exit
      -- CP-element group 21: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_Update/array_obj_ref_42_Merge/merge_req
      -- CP-element group 21: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_Update/array_obj_ref_42_Merge/merge_ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_42_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_42_load_0_ack_1, ack => accessMem_CP_0_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	1 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	24 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_48_sample_start_
      -- CP-element group 22: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_48_Sample/$entry
      -- CP-element group 22: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_48_Sample/rr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:ADD_u12_u12_48_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(22), ack => ADD_u12_u12_48_inst_req_0); -- 
    accessMem_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 14,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(24);
      gj_accessMem_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: 	32 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_48_update_start_
      -- CP-element group 23: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_48_Update/$entry
      -- CP-element group 23: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_48_Update/cr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:ADD_u12_u12_48_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(23), ack => ADD_u12_u12_48_inst_req_1); -- 
    accessMem_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(25) & accessMem_CP_0_elements(32);
      gj_accessMem_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: 	2 
    -- CP-element group 24: 	3 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_48_sample_completed_
      -- CP-element group 24: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_48_Sample/$exit
      -- CP-element group 24: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_48_Sample/ra
      -- 
    -- logger for CP element group accessMem_CP_0_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:ADD_u12_u12_48_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_48_inst_ack_0, ack => accessMem_CP_0_elements(24)); -- 
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	30 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	23 
    -- CP-element group 25:  members (29) 
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_48_update_completed_
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_48_Update/$exit
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_48_Update/ca
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_word_address_calculated
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_root_address_calculated
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_offset_calculated
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_index_resized_0
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_index_scaled_0
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_index_computed_0
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_index_resize_0/$entry
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_index_resize_0/$exit
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_index_resize_0/index_resize_req
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_index_resize_0/index_resize_ack
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_index_scale_0/$entry
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_index_scale_0/$exit
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_index_scale_0/scale_rename_req
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_index_scale_0/scale_rename_ack
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_final_index_sum_regn/$entry
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_final_index_sum_regn/$exit
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_final_index_sum_regn/req
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_final_index_sum_regn/ack
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_base_plus_offset/$entry
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_base_plus_offset/$exit
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_base_plus_offset/sum_rename_req
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_base_plus_offset/sum_rename_ack
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_word_addrgen/$entry
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_word_addrgen/$exit
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_word_addrgen/root_register_req
      -- CP-element group 25: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:ADD_u12_u12_48_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_48_inst_ack_1, ack => accessMem_CP_0_elements(25)); -- 
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	1 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	28 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_52_sample_start_
      -- CP-element group 26: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_52_Sample/$entry
      -- CP-element group 26: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_52_Sample/req
      -- 
    -- logger for CP element group accessMem_CP_0_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_47_delayed_1_0_50_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(26), ack => W_read_write_bar_47_delayed_1_0_50_inst_req_0); -- 
    accessMem_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 14,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(28);
      gj_accessMem_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: 	32 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_52_update_start_
      -- CP-element group 27: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_52_Update/$entry
      -- CP-element group 27: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_52_Update/req
      -- 
    -- logger for CP element group accessMem_CP_0_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_47_delayed_1_0_50_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(27), ack => W_read_write_bar_47_delayed_1_0_50_inst_req_1); -- 
    accessMem_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(29) & accessMem_CP_0_elements(32);
      gj_accessMem_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: 	2 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_52_sample_completed_
      -- CP-element group 28: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_52_Sample/$exit
      -- CP-element group 28: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_52_Sample/ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_47_delayed_1_0_50_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_47_delayed_1_0_50_inst_ack_0, ack => accessMem_CP_0_elements(28)); -- 
    -- CP-element group 29:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_52_update_completed_
      -- CP-element group 29: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_52_Update/$exit
      -- CP-element group 29: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_52_Update/ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_47_delayed_1_0_50_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_47_delayed_1_0_50_inst_ack_1, ack => accessMem_CP_0_elements(29)); -- 
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	25 
    -- CP-element group 30: 	29 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: 	60 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (5) 
      -- CP-element group 30: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_sample_start_
      -- CP-element group 30: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_Sample/$entry
      -- CP-element group 30: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_Sample/word_access_start/$entry
      -- CP-element group 30: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_Sample/word_access_start/word_0/$entry
      -- CP-element group 30: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_56_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(30), ack => array_obj_ref_56_load_0_req_0); -- 
    accessMem_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(25) & accessMem_CP_0_elements(29) & accessMem_CP_0_elements(32) & accessMem_CP_0_elements(60);
      gj_accessMem_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: 	56 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (5) 
      -- CP-element group 31: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_update_start_
      -- CP-element group 31: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_Update/$entry
      -- CP-element group 31: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_Update/word_access_complete/$entry
      -- CP-element group 31: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_Update/word_access_complete/word_0/$entry
      -- CP-element group 31: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_56_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(31), ack => array_obj_ref_56_load_0_req_1); -- 
    accessMem_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(33) & accessMem_CP_0_elements(56);
      gj_accessMem_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	72 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	23 
    -- CP-element group 32: 	27 
    -- CP-element group 32: 	30 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_sample_completed_
      -- CP-element group 32: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_Sample/$exit
      -- CP-element group 32: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_Sample/word_access_start/$exit
      -- CP-element group 32: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_Sample/word_access_start/word_0/$exit
      -- CP-element group 32: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group accessMem_CP_0_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_56_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_56_load_0_ack_0, ack => accessMem_CP_0_elements(32)); -- 
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	54 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (9) 
      -- CP-element group 33: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_update_completed_
      -- CP-element group 33: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_Update/$exit
      -- CP-element group 33: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_Update/word_access_complete/$exit
      -- CP-element group 33: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_Update/word_access_complete/word_0/$exit
      -- CP-element group 33: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_Update/word_access_complete/word_0/ca
      -- CP-element group 33: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_Update/array_obj_ref_56_Merge/$entry
      -- CP-element group 33: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_Update/array_obj_ref_56_Merge/$exit
      -- CP-element group 33: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_Update/array_obj_ref_56_Merge/merge_req
      -- CP-element group 33: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_Update/array_obj_ref_56_Merge/merge_ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_56_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_56_load_0_ack_1, ack => accessMem_CP_0_elements(33)); -- 
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	1 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_62_sample_start_
      -- CP-element group 34: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_62_Sample/$entry
      -- CP-element group 34: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_62_Sample/rr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:ADD_u12_u12_62_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(34), ack => ADD_u12_u12_62_inst_req_0); -- 
    accessMem_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 14,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(36);
      gj_accessMem_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	37 
    -- CP-element group 35: 	44 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_62_update_start_
      -- CP-element group 35: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_62_Update/$entry
      -- CP-element group 35: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_62_Update/cr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:ADD_u12_u12_62_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(35), ack => ADD_u12_u12_62_inst_req_1); -- 
    accessMem_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(37) & accessMem_CP_0_elements(44);
      gj_accessMem_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: 	2 
    -- CP-element group 36: 	3 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_62_sample_completed_
      -- CP-element group 36: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_62_Sample/$exit
      -- CP-element group 36: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_62_Sample/ra
      -- 
    -- logger for CP element group accessMem_CP_0_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(36) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:ADD_u12_u12_62_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_62_inst_ack_0, ack => accessMem_CP_0_elements(36)); -- 
    -- CP-element group 37:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	42 
    -- CP-element group 37: marked-successors 
    -- CP-element group 37: 	35 
    -- CP-element group 37:  members (29) 
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_index_resize_0/$entry
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_index_resize_0/$exit
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_index_resize_0/index_resize_req
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_index_resize_0/index_resize_ack
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_index_scale_0/$entry
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_index_scale_0/$exit
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_index_scale_0/scale_rename_req
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_index_scale_0/scale_rename_ack
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_final_index_sum_regn/$entry
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_final_index_sum_regn/$exit
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_final_index_sum_regn/req
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_final_index_sum_regn/ack
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_62_update_completed_
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_62_Update/$exit
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/ADD_u12_u12_62_Update/ca
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_word_address_calculated
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_root_address_calculated
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_offset_calculated
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_index_resized_0
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_index_scaled_0
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_index_computed_0
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_base_plus_offset/$entry
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_base_plus_offset/$exit
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_base_plus_offset/sum_rename_req
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_base_plus_offset/sum_rename_ack
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_word_addrgen/$entry
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_word_addrgen/$exit
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_word_addrgen/root_register_req
      -- CP-element group 37: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:ADD_u12_u12_62_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_62_inst_ack_1, ack => accessMem_CP_0_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	1 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	40 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_66_sample_start_
      -- CP-element group 38: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_66_Sample/$entry
      -- CP-element group 38: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_66_Sample/req
      -- 
    -- logger for CP element group accessMem_CP_0_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(38) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_58_delayed_1_0_64_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(38), ack => W_read_write_bar_58_delayed_1_0_64_inst_req_0); -- 
    accessMem_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 14,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(40);
      gj_accessMem_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: 	44 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_66_update_start_
      -- CP-element group 39: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_66_Update/$entry
      -- CP-element group 39: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_66_Update/req
      -- 
    -- logger for CP element group accessMem_CP_0_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_58_delayed_1_0_64_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(39), ack => W_read_write_bar_58_delayed_1_0_64_inst_req_1); -- 
    accessMem_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(41) & accessMem_CP_0_elements(44);
      gj_accessMem_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: 	2 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_66_sample_completed_
      -- CP-element group 40: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_66_Sample/$exit
      -- CP-element group 40: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_66_Sample/ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(40) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_58_delayed_1_0_64_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_58_delayed_1_0_64_inst_ack_0, ack => accessMem_CP_0_elements(40)); -- 
    -- CP-element group 41:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	39 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_66_update_completed_
      -- CP-element group 41: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_66_Update/$exit
      -- CP-element group 41: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_66_Update/ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(41) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_58_delayed_1_0_64_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_58_delayed_1_0_64_inst_ack_1, ack => accessMem_CP_0_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	37 
    -- CP-element group 42: 	41 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: 	60 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_sample_start_
      -- CP-element group 42: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_Sample/$entry
      -- CP-element group 42: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_Sample/word_access_start/$entry
      -- CP-element group 42: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_Sample/word_access_start/word_0/$entry
      -- CP-element group 42: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(42) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_70_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(42), ack => array_obj_ref_70_load_0_req_0); -- 
    accessMem_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(37) & accessMem_CP_0_elements(41) & accessMem_CP_0_elements(44) & accessMem_CP_0_elements(60);
      gj_accessMem_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	45 
    -- CP-element group 43: 	56 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (5) 
      -- CP-element group 43: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_update_start_
      -- CP-element group 43: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_Update/$entry
      -- CP-element group 43: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_Update/word_access_complete/$entry
      -- CP-element group 43: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_Update/word_access_complete/word_0/$entry
      -- CP-element group 43: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(43) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_70_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(43), ack => array_obj_ref_70_load_0_req_1); -- 
    accessMem_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(45) & accessMem_CP_0_elements(56);
      gj_accessMem_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	73 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	35 
    -- CP-element group 44: 	39 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (5) 
      -- CP-element group 44: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_sample_completed_
      -- CP-element group 44: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_Sample/$exit
      -- CP-element group 44: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_Sample/word_access_start/$exit
      -- CP-element group 44: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_Sample/word_access_start/word_0/$exit
      -- CP-element group 44: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group accessMem_CP_0_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(44) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_70_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_70_load_0_ack_0, ack => accessMem_CP_0_elements(44)); -- 
    -- CP-element group 45:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	54 
    -- CP-element group 45: marked-successors 
    -- CP-element group 45: 	43 
    -- CP-element group 45:  members (9) 
      -- CP-element group 45: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_update_completed_
      -- CP-element group 45: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_Update/$exit
      -- CP-element group 45: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_Update/word_access_complete/$exit
      -- CP-element group 45: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_Update/word_access_complete/word_0/$exit
      -- CP-element group 45: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_Update/word_access_complete/word_0/ca
      -- CP-element group 45: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_Update/array_obj_ref_70_Merge/$entry
      -- CP-element group 45: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_Update/array_obj_ref_70_Merge/$exit
      -- CP-element group 45: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_Update/array_obj_ref_70_Merge/merge_req
      -- CP-element group 45: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_Update/array_obj_ref_70_Merge/merge_ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(45) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_70_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_70_load_0_ack_1, ack => accessMem_CP_0_elements(45)); -- 
    -- CP-element group 46:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	9 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	48 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_74_sample_start_
      -- CP-element group 46: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_74_Sample/$entry
      -- CP-element group 46: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_74_Sample/req
      -- 
    -- logger for CP element group accessMem_CP_0_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(46) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_t_read_data0_69_delayed_1_0_72_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(46), ack => W_t_read_data0_69_delayed_1_0_72_inst_req_0); -- 
    accessMem_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(9) & accessMem_CP_0_elements(48);
      gj_accessMem_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	49 
    -- CP-element group 47: 	56 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_74_update_start_
      -- CP-element group 47: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_74_Update/$entry
      -- CP-element group 47: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_74_Update/req
      -- 
    -- logger for CP element group accessMem_CP_0_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(47) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_t_read_data0_69_delayed_1_0_72_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(47), ack => W_t_read_data0_69_delayed_1_0_72_inst_req_1); -- 
    accessMem_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(49) & accessMem_CP_0_elements(56);
      gj_accessMem_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: marked-successors 
    -- CP-element group 48: 	7 
    -- CP-element group 48: 	46 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_74_sample_completed_
      -- CP-element group 48: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_74_Sample/$exit
      -- CP-element group 48: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_74_Sample/ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(48) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_t_read_data0_69_delayed_1_0_72_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_t_read_data0_69_delayed_1_0_72_inst_ack_0, ack => accessMem_CP_0_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	54 
    -- CP-element group 49: marked-successors 
    -- CP-element group 49: 	47 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_74_update_completed_
      -- CP-element group 49: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_74_Update/$exit
      -- CP-element group 49: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_74_Update/ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(49) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_t_read_data0_69_delayed_1_0_72_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_t_read_data0_69_delayed_1_0_72_inst_ack_1, ack => accessMem_CP_0_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	1 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	52 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_77_sample_start_
      -- CP-element group 50: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_77_Sample/$entry
      -- CP-element group 50: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_77_Sample/req
      -- 
    -- logger for CP element group accessMem_CP_0_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(50) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_63_delayed_6_0_75_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(50), ack => W_read_write_bar_63_delayed_6_0_75_inst_req_0); -- 
    accessMem_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 14,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(52);
      gj_accessMem_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	53 
    -- CP-element group 51: 	56 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_77_update_start_
      -- CP-element group 51: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_77_Update/$entry
      -- CP-element group 51: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_77_Update/req
      -- 
    -- logger for CP element group accessMem_CP_0_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(51) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_63_delayed_6_0_75_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(51), ack => W_read_write_bar_63_delayed_6_0_75_inst_req_1); -- 
    accessMem_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(53) & accessMem_CP_0_elements(56);
      gj_accessMem_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	2 
    -- CP-element group 52: 	50 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_77_sample_completed_
      -- CP-element group 52: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_77_Sample/$exit
      -- CP-element group 52: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_77_Sample/ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(52) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_63_delayed_6_0_75_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_63_delayed_6_0_75_inst_ack_0, ack => accessMem_CP_0_elements(52)); -- 
    -- CP-element group 53:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53: marked-successors 
    -- CP-element group 53: 	51 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_77_update_completed_
      -- CP-element group 53: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_77_Update/$exit
      -- CP-element group 53: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_77_Update/ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(53) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_63_delayed_6_0_75_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_63_delayed_6_0_75_inst_ack_1, ack => accessMem_CP_0_elements(53)); -- 
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	21 
    -- CP-element group 54: 	33 
    -- CP-element group 54: 	45 
    -- CP-element group 54: 	49 
    -- CP-element group 54: 	53 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	56 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 assign_stmt_29_to_assign_stmt_101/CONCAT_u32_u64_86_sample_start_
      -- CP-element group 54: 	 assign_stmt_29_to_assign_stmt_101/CONCAT_u32_u64_86_Sample/$entry
      -- CP-element group 54: 	 assign_stmt_29_to_assign_stmt_101/CONCAT_u32_u64_86_Sample/rr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(54) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:CONCAT_u32_u64_86_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(54), ack => CONCAT_u32_u64_86_inst_req_0); -- 
    accessMem_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(21) & accessMem_CP_0_elements(33) & accessMem_CP_0_elements(45) & accessMem_CP_0_elements(49) & accessMem_CP_0_elements(53) & accessMem_CP_0_elements(56);
      gj_accessMem_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	57 
    -- CP-element group 55: 	68 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 assign_stmt_29_to_assign_stmt_101/CONCAT_u32_u64_86_update_start_
      -- CP-element group 55: 	 assign_stmt_29_to_assign_stmt_101/CONCAT_u32_u64_86_Update/$entry
      -- CP-element group 55: 	 assign_stmt_29_to_assign_stmt_101/CONCAT_u32_u64_86_Update/cr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(55) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:CONCAT_u32_u64_86_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(55), ack => CONCAT_u32_u64_86_inst_req_1); -- 
    accessMem_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(57) & accessMem_CP_0_elements(68);
      gj_accessMem_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	31 
    -- CP-element group 56: 	43 
    -- CP-element group 56: 	19 
    -- CP-element group 56: 	47 
    -- CP-element group 56: 	51 
    -- CP-element group 56: 	54 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 assign_stmt_29_to_assign_stmt_101/CONCAT_u32_u64_86_sample_completed_
      -- CP-element group 56: 	 assign_stmt_29_to_assign_stmt_101/CONCAT_u32_u64_86_Sample/$exit
      -- CP-element group 56: 	 assign_stmt_29_to_assign_stmt_101/CONCAT_u32_u64_86_Sample/ra
      -- 
    -- logger for CP element group accessMem_CP_0_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(56) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:CONCAT_u32_u64_86_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_86_inst_ack_0, ack => accessMem_CP_0_elements(56)); -- 
    -- CP-element group 57:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	66 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	55 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 assign_stmt_29_to_assign_stmt_101/CONCAT_u32_u64_86_update_completed_
      -- CP-element group 57: 	 assign_stmt_29_to_assign_stmt_101/CONCAT_u32_u64_86_Update/$exit
      -- CP-element group 57: 	 assign_stmt_29_to_assign_stmt_101/CONCAT_u32_u64_86_Update/ca
      -- 
    -- logger for CP element group accessMem_CP_0_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(57) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:CONCAT_u32_u64_86_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_86_inst_ack_1, ack => accessMem_CP_0_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	1 
    -- CP-element group 58: 	70 
    -- CP-element group 58: 	71 
    -- CP-element group 58: 	72 
    -- CP-element group 58: 	73 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_sample_start_
      -- CP-element group 58: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_Sample/$entry
      -- CP-element group 58: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_Sample/array_obj_ref_90_Split/$entry
      -- CP-element group 58: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_Sample/array_obj_ref_90_Split/$exit
      -- CP-element group 58: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_Sample/array_obj_ref_90_Split/split_req
      -- CP-element group 58: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_Sample/array_obj_ref_90_Split/split_ack
      -- CP-element group 58: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_Sample/word_access_start/$entry
      -- CP-element group 58: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_Sample/word_access_start/word_0/$entry
      -- CP-element group 58: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(58) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_90_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(58), ack => array_obj_ref_90_store_0_req_0); -- 
    accessMem_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 14,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(70) & accessMem_CP_0_elements(71) & accessMem_CP_0_elements(72) & accessMem_CP_0_elements(73) & accessMem_CP_0_elements(60);
      gj_accessMem_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (5) 
      -- CP-element group 59: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_update_start_
      -- CP-element group 59: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_Update/$entry
      -- CP-element group 59: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_Update/word_access_complete/$entry
      -- CP-element group 59: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_Update/word_access_complete/word_0/$entry
      -- CP-element group 59: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(59) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_90_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(59), ack => array_obj_ref_90_store_0_req_1); -- 
    accessMem_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMem_CP_0_elements(61);
      gj_accessMem_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	74 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	30 
    -- CP-element group 60: 	42 
    -- CP-element group 60: 	2 
    -- CP-element group 60: 	3 
    -- CP-element group 60: 	4 
    -- CP-element group 60: 	6 
    -- CP-element group 60: 	18 
    -- CP-element group 60: 	58 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_sample_completed_
      -- CP-element group 60: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_Sample/$exit
      -- CP-element group 60: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_Sample/word_access_start/$exit
      -- CP-element group 60: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_Sample/word_access_start/word_0/$exit
      -- CP-element group 60: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_Sample/word_access_start/word_0/ra
      -- CP-element group 60: 	 assign_stmt_29_to_assign_stmt_101/ring_reenable_memory_space_5
      -- 
    -- logger for CP element group accessMem_CP_0_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(60) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_90_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_90_store_0_ack_0, ack => accessMem_CP_0_elements(60)); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	74 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (5) 
      -- CP-element group 61: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_update_completed_
      -- CP-element group 61: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_Update/$exit
      -- CP-element group 61: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_Update/word_access_complete/$exit
      -- CP-element group 61: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_Update/word_access_complete/word_0/$exit
      -- CP-element group 61: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_90_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group accessMem_CP_0_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(61) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_90_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_90_store_0_ack_1, ack => accessMem_CP_0_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	1 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_95_sample_start_
      -- CP-element group 62: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_95_Sample/$entry
      -- CP-element group 62: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_95_Sample/req
      -- 
    -- logger for CP element group accessMem_CP_0_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(62) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_79_delayed_7_0_93_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(62), ack => W_read_write_bar_79_delayed_7_0_93_inst_req_0); -- 
    accessMem_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 14,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(64);
      gj_accessMem_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: 	68 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_95_update_start_
      -- CP-element group 63: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_95_Update/$entry
      -- CP-element group 63: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_95_Update/req
      -- 
    -- logger for CP element group accessMem_CP_0_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(63) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_79_delayed_7_0_93_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(63), ack => W_read_write_bar_79_delayed_7_0_93_inst_req_1); -- 
    accessMem_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(65) & accessMem_CP_0_elements(68);
      gj_accessMem_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	2 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_95_sample_completed_
      -- CP-element group 64: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_95_Sample/$exit
      -- CP-element group 64: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_95_Sample/ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(64) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_79_delayed_7_0_93_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_79_delayed_7_0_93_inst_ack_0, ack => accessMem_CP_0_elements(64)); -- 
    -- CP-element group 65:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65: marked-successors 
    -- CP-element group 65: 	63 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_95_update_completed_
      -- CP-element group 65: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_95_Update/$exit
      -- CP-element group 65: 	 assign_stmt_29_to_assign_stmt_101/assign_stmt_95_Update/ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(65) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_79_delayed_7_0_93_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_79_delayed_7_0_93_inst_ack_1, ack => accessMem_CP_0_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	57 
    -- CP-element group 66: 	65 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	68 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 assign_stmt_29_to_assign_stmt_101/MUX_100_sample_start_
      -- CP-element group 66: 	 assign_stmt_29_to_assign_stmt_101/MUX_100_start/$entry
      -- CP-element group 66: 	 assign_stmt_29_to_assign_stmt_101/MUX_100_start/req
      -- 
    -- logger for CP element group accessMem_CP_0_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(66) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:MUX_100_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(66), ack => MUX_100_inst_req_0); -- 
    accessMem_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(57) & accessMem_CP_0_elements(65) & accessMem_CP_0_elements(68);
      gj_accessMem_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	5 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 assign_stmt_29_to_assign_stmt_101/MUX_100_update_start_
      -- CP-element group 67: 	 assign_stmt_29_to_assign_stmt_101/MUX_100_complete/$entry
      -- CP-element group 67: 	 assign_stmt_29_to_assign_stmt_101/MUX_100_complete/req
      -- 
    -- logger for CP element group accessMem_CP_0_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(67) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:MUX_100_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(67), ack => MUX_100_inst_req_1); -- 
    accessMem_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 14,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(5) & accessMem_CP_0_elements(69);
      gj_accessMem_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	55 
    -- CP-element group 68: 	63 
    -- CP-element group 68: 	66 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 assign_stmt_29_to_assign_stmt_101/MUX_100_sample_completed_
      -- CP-element group 68: 	 assign_stmt_29_to_assign_stmt_101/MUX_100_start/$exit
      -- CP-element group 68: 	 assign_stmt_29_to_assign_stmt_101/MUX_100_start/ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(68) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:MUX_100_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_100_inst_ack_0, ack => accessMem_CP_0_elements(68)); -- 
    -- CP-element group 69:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	74 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	67 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 assign_stmt_29_to_assign_stmt_101/MUX_100_update_completed_
      -- CP-element group 69: 	 assign_stmt_29_to_assign_stmt_101/MUX_100_complete/$exit
      -- CP-element group 69: 	 assign_stmt_29_to_assign_stmt_101/MUX_100_complete/ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(69) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:MUX_100_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_100_inst_ack_1, ack => accessMem_CP_0_elements(69)); -- 
    -- CP-element group 70:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	8 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	58 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_28_array_obj_ref_90_delay
      -- 
    -- logger for CP element group accessMem_CP_0_elements(70)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(70)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(70) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accessMem_CP_0_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => accessMem_CP_0_elements(8), ack => accessMem_CP_0_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	20 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	58 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_42_array_obj_ref_90_delay
      -- 
    -- logger for CP element group accessMem_CP_0_elements(71)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(71)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(71) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accessMem_CP_0_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => accessMem_CP_0_elements(20), ack => accessMem_CP_0_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	32 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	58 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_56_array_obj_ref_90_delay
      -- 
    -- logger for CP element group accessMem_CP_0_elements(72)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(72)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(72) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accessMem_CP_0_elements(72) is a control-delay.
    cp_element_72_delay: control_delay_element  generic map(name => " 72_delay", delay_value => 1)  port map(req => accessMem_CP_0_elements(32), ack => accessMem_CP_0_elements(72), clk => clk, reset =>reset);
    -- CP-element group 73:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	44 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	58 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 assign_stmt_29_to_assign_stmt_101/array_obj_ref_70_array_obj_ref_90_delay
      -- 
    -- logger for CP element group accessMem_CP_0_elements(73)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(73)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(73) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accessMem_CP_0_elements(73) is a control-delay.
    cp_element_73_delay: control_delay_element  generic map(name => " 73_delay", delay_value => 1)  port map(req => accessMem_CP_0_elements(44), ack => accessMem_CP_0_elements(73), clk => clk, reset =>reset);
    -- CP-element group 74:  join  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	60 
    -- CP-element group 74: 	61 
    -- CP-element group 74: 	69 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	79 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 assign_stmt_29_to_assign_stmt_101/$exit
      -- 
    -- logger for CP element group accessMem_CP_0_elements(74)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(74)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(74) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 14,1 => 14,2 => 14);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(60) & accessMem_CP_0_elements(61) & accessMem_CP_0_elements(69);
      gj_accessMem_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  place  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	2 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 read_write_bar_update_enable
      -- 
    -- logger for CP element group accessMem_CP_0_elements(75)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(75)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(75) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_CP_0_elements(75) <= accessMem_CP_0_elements(2);
    -- CP-element group 76:  place  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	3 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 addr_update_enable
      -- 
    -- logger for CP element group accessMem_CP_0_elements(76)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(76)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(76) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_CP_0_elements(76) <= accessMem_CP_0_elements(3);
    -- CP-element group 77:  place  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	4 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 write_data_update_enable
      -- 
    -- logger for CP element group accessMem_CP_0_elements(77)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(77)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(77) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_CP_0_elements(77) <= accessMem_CP_0_elements(4);
    -- CP-element group 78:  place  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	5 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 read_datal_update_enable
      -- 
    -- logger for CP element group accessMem_CP_0_elements(78)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(78)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(78) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 79:  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	74 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 $exit
      -- 
    -- logger for CP element group accessMem_CP_0_elements(79)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(79)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(79) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_CP_0_elements(79) <= accessMem_CP_0_elements(74);
    --  hookup: inputs to control-path 
    accessMem_CP_0_elements(78) <= read_datal_update_enable;
    -- hookup: output from control-path 
    read_write_bar_update_enable <= accessMem_CP_0_elements(75);
    addr_update_enable <= accessMem_CP_0_elements(76);
    write_data_update_enable <= accessMem_CP_0_elements(77);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u16_u32_82_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_85_wire : std_logic_vector(31 downto 0);
    signal R_addr1_41_resized : std_logic_vector(10 downto 0);
    signal R_addr1_41_scaled : std_logic_vector(10 downto 0);
    signal R_addr2_55_resized : std_logic_vector(10 downto 0);
    signal R_addr2_55_scaled : std_logic_vector(10 downto 0);
    signal R_addr3_69_resized : std_logic_vector(10 downto 0);
    signal R_addr3_69_scaled : std_logic_vector(10 downto 0);
    signal R_addr_27_resized : std_logic_vector(10 downto 0);
    signal R_addr_27_scaled : std_logic_vector(10 downto 0);
    signal R_addr_89_resized : std_logic_vector(10 downto 0);
    signal R_addr_89_scaled : std_logic_vector(10 downto 0);
    signal addr1_35 : std_logic_vector(11 downto 0);
    signal addr2_49 : std_logic_vector(11 downto 0);
    signal addr3_63 : std_logic_vector(11 downto 0);
    signal array_obj_ref_28_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_28_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_28_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_28_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_28_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_28_word_address_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_28_word_offset_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_42_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_42_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_42_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_42_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_42_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_42_word_address_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_42_word_offset_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_56_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_56_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_56_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_56_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_56_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_56_word_address_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_56_word_offset_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_70_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_70_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_70_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_70_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_70_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_70_word_address_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_70_word_offset_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_90_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_90_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_90_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_90_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_90_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_90_word_address_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_90_word_offset_0 : std_logic_vector(10 downto 0);
    signal konst_33_wire_constant : std_logic_vector(11 downto 0);
    signal konst_47_wire_constant : std_logic_vector(11 downto 0);
    signal konst_61_wire_constant : std_logic_vector(11 downto 0);
    signal konst_99_wire_constant : std_logic_vector(63 downto 0);
    signal read_write_bar_36_delayed_1_0_38 : std_logic_vector(0 downto 0);
    signal read_write_bar_47_delayed_1_0_52 : std_logic_vector(0 downto 0);
    signal read_write_bar_58_delayed_1_0_66 : std_logic_vector(0 downto 0);
    signal read_write_bar_63_delayed_6_0_77 : std_logic_vector(0 downto 0);
    signal read_write_bar_79_delayed_7_0_95 : std_logic_vector(0 downto 0);
    signal t_read_data0_29 : std_logic_vector(15 downto 0);
    signal t_read_data0_69_delayed_1_0_74 : std_logic_vector(15 downto 0);
    signal t_read_data1_43 : std_logic_vector(15 downto 0);
    signal t_read_data2_57 : std_logic_vector(15 downto 0);
    signal t_read_data3_71 : std_logic_vector(15 downto 0);
    signal t_read_datal_87 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_28_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_28_resized_base_address <= "00000000000";
    array_obj_ref_28_word_offset_0 <= "00000000000";
    array_obj_ref_42_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_42_resized_base_address <= "00000000000";
    array_obj_ref_42_word_offset_0 <= "00000000000";
    array_obj_ref_56_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_56_resized_base_address <= "00000000000";
    array_obj_ref_56_word_offset_0 <= "00000000000";
    array_obj_ref_70_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_70_resized_base_address <= "00000000000";
    array_obj_ref_70_word_offset_0 <= "00000000000";
    array_obj_ref_90_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_90_resized_base_address <= "00000000000";
    array_obj_ref_90_word_offset_0 <= "00000000000";
    konst_33_wire_constant <= "000000000001";
    konst_47_wire_constant <= "000000000010";
    konst_61_wire_constant <= "000000000011";
    konst_99_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- logger for split-operator MUX_100_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if MUX_100_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:MUX_100_inst:started:   inputs: " & " read_write_bar_79_delayed_7_0_95 = "& Convert_SLV_To_Hex_String(read_write_bar_79_delayed_7_0_95) & " t_read_datal_87 = "& Convert_SLV_To_Hex_String(t_read_datal_87) & " konst_99_wire_constant = "& Convert_SLV_To_Hex_String(konst_99_wire_constant));
          --
        end if; 
        if MUX_100_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:MUX_100_inst:finished:  outputs: " & " read_datal_buffer= "  & Convert_SLV_To_Hex_String(read_datal_buffer));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    MUX_100_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_100_inst_req_0;
      MUX_100_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_100_inst_req_1;
      MUX_100_inst_ack_1<= update_ack(0);
      MUX_100_inst: SelectSplitProtocol generic map(name => "MUX_100_inst", data_width => 64, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => t_read_datal_87, y => konst_99_wire_constant, sel => read_write_bar_79_delayed_7_0_95, z => read_datal_buffer, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator W_read_write_bar_36_delayed_1_0_36_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_read_write_bar_36_delayed_1_0_36_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:W_read_write_bar_36_delayed_1_0_36_inst:started:   inputs: " & " read_write_bar_buffer = "& Convert_SLV_To_Hex_String(read_write_bar_buffer));
          --
        end if; 
        if W_read_write_bar_36_delayed_1_0_36_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:W_read_write_bar_36_delayed_1_0_36_inst:finished:  outputs: " & " read_write_bar_36_delayed_1_0_38= "  & Convert_SLV_To_Hex_String(read_write_bar_36_delayed_1_0_38));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_read_write_bar_36_delayed_1_0_36_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_write_bar_36_delayed_1_0_36_inst_req_0;
      W_read_write_bar_36_delayed_1_0_36_inst_ack_0<= wack(0);
      rreq(0) <= W_read_write_bar_36_delayed_1_0_36_inst_req_1;
      W_read_write_bar_36_delayed_1_0_36_inst_ack_1<= rack(0);
      W_read_write_bar_36_delayed_1_0_36_inst : InterlockBuffer generic map ( -- 
        name => "W_read_write_bar_36_delayed_1_0_36_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_write_bar_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_write_bar_36_delayed_1_0_38,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_read_write_bar_47_delayed_1_0_50_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_read_write_bar_47_delayed_1_0_50_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:W_read_write_bar_47_delayed_1_0_50_inst:started:   inputs: " & " read_write_bar_buffer = "& Convert_SLV_To_Hex_String(read_write_bar_buffer));
          --
        end if; 
        if W_read_write_bar_47_delayed_1_0_50_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:W_read_write_bar_47_delayed_1_0_50_inst:finished:  outputs: " & " read_write_bar_47_delayed_1_0_52= "  & Convert_SLV_To_Hex_String(read_write_bar_47_delayed_1_0_52));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_read_write_bar_47_delayed_1_0_50_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_write_bar_47_delayed_1_0_50_inst_req_0;
      W_read_write_bar_47_delayed_1_0_50_inst_ack_0<= wack(0);
      rreq(0) <= W_read_write_bar_47_delayed_1_0_50_inst_req_1;
      W_read_write_bar_47_delayed_1_0_50_inst_ack_1<= rack(0);
      W_read_write_bar_47_delayed_1_0_50_inst : InterlockBuffer generic map ( -- 
        name => "W_read_write_bar_47_delayed_1_0_50_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_write_bar_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_write_bar_47_delayed_1_0_52,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_read_write_bar_58_delayed_1_0_64_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_read_write_bar_58_delayed_1_0_64_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:W_read_write_bar_58_delayed_1_0_64_inst:started:   inputs: " & " read_write_bar_buffer = "& Convert_SLV_To_Hex_String(read_write_bar_buffer));
          --
        end if; 
        if W_read_write_bar_58_delayed_1_0_64_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:W_read_write_bar_58_delayed_1_0_64_inst:finished:  outputs: " & " read_write_bar_58_delayed_1_0_66= "  & Convert_SLV_To_Hex_String(read_write_bar_58_delayed_1_0_66));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_read_write_bar_58_delayed_1_0_64_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_write_bar_58_delayed_1_0_64_inst_req_0;
      W_read_write_bar_58_delayed_1_0_64_inst_ack_0<= wack(0);
      rreq(0) <= W_read_write_bar_58_delayed_1_0_64_inst_req_1;
      W_read_write_bar_58_delayed_1_0_64_inst_ack_1<= rack(0);
      W_read_write_bar_58_delayed_1_0_64_inst : InterlockBuffer generic map ( -- 
        name => "W_read_write_bar_58_delayed_1_0_64_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_write_bar_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_write_bar_58_delayed_1_0_66,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_read_write_bar_63_delayed_6_0_75_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_read_write_bar_63_delayed_6_0_75_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:W_read_write_bar_63_delayed_6_0_75_inst:started:   inputs: " & " read_write_bar_buffer = "& Convert_SLV_To_Hex_String(read_write_bar_buffer));
          --
        end if; 
        if W_read_write_bar_63_delayed_6_0_75_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:W_read_write_bar_63_delayed_6_0_75_inst:finished:  outputs: " & " read_write_bar_63_delayed_6_0_77= "  & Convert_SLV_To_Hex_String(read_write_bar_63_delayed_6_0_77));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_read_write_bar_63_delayed_6_0_75_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_write_bar_63_delayed_6_0_75_inst_req_0;
      W_read_write_bar_63_delayed_6_0_75_inst_ack_0<= wack(0);
      rreq(0) <= W_read_write_bar_63_delayed_6_0_75_inst_req_1;
      W_read_write_bar_63_delayed_6_0_75_inst_ack_1<= rack(0);
      W_read_write_bar_63_delayed_6_0_75_inst : InterlockBuffer generic map ( -- 
        name => "W_read_write_bar_63_delayed_6_0_75_inst",
        buffer_size => 6,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_write_bar_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_write_bar_63_delayed_6_0_77,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_read_write_bar_79_delayed_7_0_93_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_read_write_bar_79_delayed_7_0_93_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:W_read_write_bar_79_delayed_7_0_93_inst:started:   inputs: " & " read_write_bar_buffer = "& Convert_SLV_To_Hex_String(read_write_bar_buffer));
          --
        end if; 
        if W_read_write_bar_79_delayed_7_0_93_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:W_read_write_bar_79_delayed_7_0_93_inst:finished:  outputs: " & " read_write_bar_79_delayed_7_0_95= "  & Convert_SLV_To_Hex_String(read_write_bar_79_delayed_7_0_95));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_read_write_bar_79_delayed_7_0_93_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_write_bar_79_delayed_7_0_93_inst_req_0;
      W_read_write_bar_79_delayed_7_0_93_inst_ack_0<= wack(0);
      rreq(0) <= W_read_write_bar_79_delayed_7_0_93_inst_req_1;
      W_read_write_bar_79_delayed_7_0_93_inst_ack_1<= rack(0);
      W_read_write_bar_79_delayed_7_0_93_inst : InterlockBuffer generic map ( -- 
        name => "W_read_write_bar_79_delayed_7_0_93_inst",
        buffer_size => 7,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_write_bar_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_write_bar_79_delayed_7_0_95,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_t_read_data0_69_delayed_1_0_72_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_t_read_data0_69_delayed_1_0_72_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:W_t_read_data0_69_delayed_1_0_72_inst:started:   inputs: " & " t_read_data0_29 = "& Convert_SLV_To_Hex_String(t_read_data0_29));
          --
        end if; 
        if W_t_read_data0_69_delayed_1_0_72_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:W_t_read_data0_69_delayed_1_0_72_inst:finished:  outputs: " & " t_read_data0_69_delayed_1_0_74= "  & Convert_SLV_To_Hex_String(t_read_data0_69_delayed_1_0_74));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_t_read_data0_69_delayed_1_0_72_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_t_read_data0_69_delayed_1_0_72_inst_req_0;
      W_t_read_data0_69_delayed_1_0_72_inst_ack_0<= wack(0);
      rreq(0) <= W_t_read_data0_69_delayed_1_0_72_inst_req_1;
      W_t_read_data0_69_delayed_1_0_72_inst_ack_1<= rack(0);
      W_t_read_data0_69_delayed_1_0_72_inst : InterlockBuffer generic map ( -- 
        name => "W_t_read_data0_69_delayed_1_0_72_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => t_read_data0_29,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => t_read_data0_69_delayed_1_0_74,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for operator array_obj_ref_28_addr_0 flow-through 
    process(array_obj_ref_28_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_28_addr_0:flowthrough  inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " array_obj_ref_28_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_28_root_address) & "outputs: " & " array_obj_ref_28_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_28_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_28_addr_0
    process(array_obj_ref_28_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_28_root_address;
      ov(10 downto 0) := iv;
      array_obj_ref_28_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_28_gather_scatter flow-through 
    process(t_read_data0_29) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_28_gather_scatter:flowthrough  inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " array_obj_ref_28_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_28_data_0) & "outputs: " & " t_read_data0_29= "  & Convert_SLV_To_Hex_String(t_read_data0_29));
      --
    end process; 
    -- equivalence array_obj_ref_28_gather_scatter
    process(array_obj_ref_28_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_28_data_0;
      ov(15 downto 0) := iv;
      t_read_data0_29 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_28_index_0_rename flow-through 
    process(R_addr_27_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_28_index_0_rename:flowthrough  inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " R_addr_27_resized = "& Convert_SLV_To_Hex_String(R_addr_27_resized) & "outputs: " & " R_addr_27_scaled= "  & Convert_SLV_To_Hex_String(R_addr_27_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_28_index_0_rename
    process(R_addr_27_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_27_resized;
      ov(10 downto 0) := iv;
      R_addr_27_scaled <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_28_index_0_resize flow-through 
    process(R_addr_27_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_28_index_0_resize:flowthrough  inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " addr_buffer = "& Convert_SLV_To_Hex_String(addr_buffer) & "outputs: " & " R_addr_27_resized= "  & Convert_SLV_To_Hex_String(R_addr_27_resized));
      --
    end process; 
    -- equivalence array_obj_ref_28_index_0_resize
    process(addr_buffer) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_buffer;
      ov := iv(10 downto 0);
      R_addr_27_resized <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_28_index_offset flow-through 
    process(array_obj_ref_28_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_28_index_offset:flowthrough  inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " R_addr_27_scaled = "& Convert_SLV_To_Hex_String(R_addr_27_scaled) & "outputs: " & " array_obj_ref_28_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_28_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_28_index_offset
    process(R_addr_27_scaled) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_27_scaled;
      ov(10 downto 0) := iv;
      array_obj_ref_28_final_offset <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_28_root_address_inst flow-through 
    process(array_obj_ref_28_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_28_root_address_inst:flowthrough  inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " array_obj_ref_28_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_28_final_offset) & "outputs: " & " array_obj_ref_28_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_28_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_28_root_address_inst
    process(array_obj_ref_28_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_28_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_28_root_address <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_42_addr_0 flow-through 
    process(array_obj_ref_42_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_42_addr_0:flowthrough  inputs: " & " read_write_bar_36_delayed_1_0_38 (guard)= " & Convert_SLV_To_String(read_write_bar_36_delayed_1_0_38) & " array_obj_ref_42_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_42_root_address) & "outputs: " & " array_obj_ref_42_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_42_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_42_addr_0
    process(array_obj_ref_42_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_42_root_address;
      ov(10 downto 0) := iv;
      array_obj_ref_42_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_42_gather_scatter flow-through 
    process(t_read_data1_43) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_42_gather_scatter:flowthrough  inputs: " & " read_write_bar_36_delayed_1_0_38 (guard)= " & Convert_SLV_To_String(read_write_bar_36_delayed_1_0_38) & " array_obj_ref_42_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_42_data_0) & "outputs: " & " t_read_data1_43= "  & Convert_SLV_To_Hex_String(t_read_data1_43));
      --
    end process; 
    -- equivalence array_obj_ref_42_gather_scatter
    process(array_obj_ref_42_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_42_data_0;
      ov(15 downto 0) := iv;
      t_read_data1_43 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_42_index_0_rename flow-through 
    process(R_addr1_41_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_42_index_0_rename:flowthrough  inputs: " & " read_write_bar_36_delayed_1_0_38 (guard)= " & Convert_SLV_To_String(read_write_bar_36_delayed_1_0_38) & " R_addr1_41_resized = "& Convert_SLV_To_Hex_String(R_addr1_41_resized) & "outputs: " & " R_addr1_41_scaled= "  & Convert_SLV_To_Hex_String(R_addr1_41_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_42_index_0_rename
    process(R_addr1_41_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr1_41_resized;
      ov(10 downto 0) := iv;
      R_addr1_41_scaled <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_42_index_0_resize flow-through 
    process(R_addr1_41_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_42_index_0_resize:flowthrough  inputs: " & " read_write_bar_36_delayed_1_0_38 (guard)= " & Convert_SLV_To_String(read_write_bar_36_delayed_1_0_38) & " addr1_35 = "& Convert_SLV_To_Hex_String(addr1_35) & "outputs: " & " R_addr1_41_resized= "  & Convert_SLV_To_Hex_String(R_addr1_41_resized));
      --
    end process; 
    -- equivalence array_obj_ref_42_index_0_resize
    process(addr1_35) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr1_35;
      ov := iv(10 downto 0);
      R_addr1_41_resized <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_42_index_offset flow-through 
    process(array_obj_ref_42_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_42_index_offset:flowthrough  inputs: " & " read_write_bar_36_delayed_1_0_38 (guard)= " & Convert_SLV_To_String(read_write_bar_36_delayed_1_0_38) & " R_addr1_41_scaled = "& Convert_SLV_To_Hex_String(R_addr1_41_scaled) & "outputs: " & " array_obj_ref_42_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_42_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_42_index_offset
    process(R_addr1_41_scaled) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr1_41_scaled;
      ov(10 downto 0) := iv;
      array_obj_ref_42_final_offset <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_42_root_address_inst flow-through 
    process(array_obj_ref_42_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_42_root_address_inst:flowthrough  inputs: " & " read_write_bar_36_delayed_1_0_38 (guard)= " & Convert_SLV_To_String(read_write_bar_36_delayed_1_0_38) & " array_obj_ref_42_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_42_final_offset) & "outputs: " & " array_obj_ref_42_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_42_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_42_root_address_inst
    process(array_obj_ref_42_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_42_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_42_root_address <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_56_addr_0 flow-through 
    process(array_obj_ref_56_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_56_addr_0:flowthrough  inputs: " & " read_write_bar_47_delayed_1_0_52 (guard)= " & Convert_SLV_To_String(read_write_bar_47_delayed_1_0_52) & " array_obj_ref_56_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_56_root_address) & "outputs: " & " array_obj_ref_56_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_56_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_56_addr_0
    process(array_obj_ref_56_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_56_root_address;
      ov(10 downto 0) := iv;
      array_obj_ref_56_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_56_gather_scatter flow-through 
    process(t_read_data2_57) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_56_gather_scatter:flowthrough  inputs: " & " read_write_bar_47_delayed_1_0_52 (guard)= " & Convert_SLV_To_String(read_write_bar_47_delayed_1_0_52) & " array_obj_ref_56_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_56_data_0) & "outputs: " & " t_read_data2_57= "  & Convert_SLV_To_Hex_String(t_read_data2_57));
      --
    end process; 
    -- equivalence array_obj_ref_56_gather_scatter
    process(array_obj_ref_56_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_56_data_0;
      ov(15 downto 0) := iv;
      t_read_data2_57 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_56_index_0_rename flow-through 
    process(R_addr2_55_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_56_index_0_rename:flowthrough  inputs: " & " read_write_bar_47_delayed_1_0_52 (guard)= " & Convert_SLV_To_String(read_write_bar_47_delayed_1_0_52) & " R_addr2_55_resized = "& Convert_SLV_To_Hex_String(R_addr2_55_resized) & "outputs: " & " R_addr2_55_scaled= "  & Convert_SLV_To_Hex_String(R_addr2_55_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_56_index_0_rename
    process(R_addr2_55_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr2_55_resized;
      ov(10 downto 0) := iv;
      R_addr2_55_scaled <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_56_index_0_resize flow-through 
    process(R_addr2_55_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_56_index_0_resize:flowthrough  inputs: " & " read_write_bar_47_delayed_1_0_52 (guard)= " & Convert_SLV_To_String(read_write_bar_47_delayed_1_0_52) & " addr2_49 = "& Convert_SLV_To_Hex_String(addr2_49) & "outputs: " & " R_addr2_55_resized= "  & Convert_SLV_To_Hex_String(R_addr2_55_resized));
      --
    end process; 
    -- equivalence array_obj_ref_56_index_0_resize
    process(addr2_49) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr2_49;
      ov := iv(10 downto 0);
      R_addr2_55_resized <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_56_index_offset flow-through 
    process(array_obj_ref_56_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_56_index_offset:flowthrough  inputs: " & " read_write_bar_47_delayed_1_0_52 (guard)= " & Convert_SLV_To_String(read_write_bar_47_delayed_1_0_52) & " R_addr2_55_scaled = "& Convert_SLV_To_Hex_String(R_addr2_55_scaled) & "outputs: " & " array_obj_ref_56_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_56_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_56_index_offset
    process(R_addr2_55_scaled) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr2_55_scaled;
      ov(10 downto 0) := iv;
      array_obj_ref_56_final_offset <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_56_root_address_inst flow-through 
    process(array_obj_ref_56_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_56_root_address_inst:flowthrough  inputs: " & " read_write_bar_47_delayed_1_0_52 (guard)= " & Convert_SLV_To_String(read_write_bar_47_delayed_1_0_52) & " array_obj_ref_56_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_56_final_offset) & "outputs: " & " array_obj_ref_56_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_56_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_56_root_address_inst
    process(array_obj_ref_56_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_56_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_56_root_address <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_70_addr_0 flow-through 
    process(array_obj_ref_70_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_70_addr_0:flowthrough  inputs: " & " read_write_bar_58_delayed_1_0_66 (guard)= " & Convert_SLV_To_String(read_write_bar_58_delayed_1_0_66) & " array_obj_ref_70_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_70_root_address) & "outputs: " & " array_obj_ref_70_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_70_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_70_addr_0
    process(array_obj_ref_70_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_70_root_address;
      ov(10 downto 0) := iv;
      array_obj_ref_70_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_70_gather_scatter flow-through 
    process(t_read_data3_71) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_70_gather_scatter:flowthrough  inputs: " & " read_write_bar_58_delayed_1_0_66 (guard)= " & Convert_SLV_To_String(read_write_bar_58_delayed_1_0_66) & " array_obj_ref_70_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_70_data_0) & "outputs: " & " t_read_data3_71= "  & Convert_SLV_To_Hex_String(t_read_data3_71));
      --
    end process; 
    -- equivalence array_obj_ref_70_gather_scatter
    process(array_obj_ref_70_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_70_data_0;
      ov(15 downto 0) := iv;
      t_read_data3_71 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_70_index_0_rename flow-through 
    process(R_addr3_69_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_70_index_0_rename:flowthrough  inputs: " & " read_write_bar_58_delayed_1_0_66 (guard)= " & Convert_SLV_To_String(read_write_bar_58_delayed_1_0_66) & " R_addr3_69_resized = "& Convert_SLV_To_Hex_String(R_addr3_69_resized) & "outputs: " & " R_addr3_69_scaled= "  & Convert_SLV_To_Hex_String(R_addr3_69_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_70_index_0_rename
    process(R_addr3_69_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr3_69_resized;
      ov(10 downto 0) := iv;
      R_addr3_69_scaled <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_70_index_0_resize flow-through 
    process(R_addr3_69_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_70_index_0_resize:flowthrough  inputs: " & " read_write_bar_58_delayed_1_0_66 (guard)= " & Convert_SLV_To_String(read_write_bar_58_delayed_1_0_66) & " addr3_63 = "& Convert_SLV_To_Hex_String(addr3_63) & "outputs: " & " R_addr3_69_resized= "  & Convert_SLV_To_Hex_String(R_addr3_69_resized));
      --
    end process; 
    -- equivalence array_obj_ref_70_index_0_resize
    process(addr3_63) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr3_63;
      ov := iv(10 downto 0);
      R_addr3_69_resized <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_70_index_offset flow-through 
    process(array_obj_ref_70_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_70_index_offset:flowthrough  inputs: " & " read_write_bar_58_delayed_1_0_66 (guard)= " & Convert_SLV_To_String(read_write_bar_58_delayed_1_0_66) & " R_addr3_69_scaled = "& Convert_SLV_To_Hex_String(R_addr3_69_scaled) & "outputs: " & " array_obj_ref_70_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_70_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_70_index_offset
    process(R_addr3_69_scaled) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr3_69_scaled;
      ov(10 downto 0) := iv;
      array_obj_ref_70_final_offset <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_70_root_address_inst flow-through 
    process(array_obj_ref_70_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_70_root_address_inst:flowthrough  inputs: " & " read_write_bar_58_delayed_1_0_66 (guard)= " & Convert_SLV_To_String(read_write_bar_58_delayed_1_0_66) & " array_obj_ref_70_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_70_final_offset) & "outputs: " & " array_obj_ref_70_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_70_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_70_root_address_inst
    process(array_obj_ref_70_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_70_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_70_root_address <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_90_addr_0 flow-through 
    process(array_obj_ref_90_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_90_addr_0:flowthrough  inputs: " & " read_write_bar_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_buffer) & " array_obj_ref_90_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_90_root_address) & "outputs: " & " array_obj_ref_90_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_90_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_90_addr_0
    process(array_obj_ref_90_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_90_root_address;
      ov(10 downto 0) := iv;
      array_obj_ref_90_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_90_gather_scatter flow-through 
    process(array_obj_ref_90_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_90_gather_scatter:flowthrough  inputs: " & " read_write_bar_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_buffer) & " write_data_buffer = "& Convert_SLV_To_Hex_String(write_data_buffer) & "outputs: " & " array_obj_ref_90_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_90_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_90_gather_scatter
    process(write_data_buffer) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := write_data_buffer;
      ov(15 downto 0) := iv;
      array_obj_ref_90_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_90_index_0_rename flow-through 
    process(R_addr_89_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_90_index_0_rename:flowthrough  inputs: " & " read_write_bar_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_buffer) & " R_addr_89_resized = "& Convert_SLV_To_Hex_String(R_addr_89_resized) & "outputs: " & " R_addr_89_scaled= "  & Convert_SLV_To_Hex_String(R_addr_89_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_90_index_0_rename
    process(R_addr_89_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_89_resized;
      ov(10 downto 0) := iv;
      R_addr_89_scaled <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_90_index_0_resize flow-through 
    process(R_addr_89_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_90_index_0_resize:flowthrough  inputs: " & " read_write_bar_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_buffer) & " addr_buffer = "& Convert_SLV_To_Hex_String(addr_buffer) & "outputs: " & " R_addr_89_resized= "  & Convert_SLV_To_Hex_String(R_addr_89_resized));
      --
    end process; 
    -- equivalence array_obj_ref_90_index_0_resize
    process(addr_buffer) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_buffer;
      ov := iv(10 downto 0);
      R_addr_89_resized <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_90_index_offset flow-through 
    process(array_obj_ref_90_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_90_index_offset:flowthrough  inputs: " & " read_write_bar_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_buffer) & " R_addr_89_scaled = "& Convert_SLV_To_Hex_String(R_addr_89_scaled) & "outputs: " & " array_obj_ref_90_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_90_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_90_index_offset
    process(R_addr_89_scaled) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_89_scaled;
      ov(10 downto 0) := iv;
      array_obj_ref_90_final_offset <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_90_root_address_inst flow-through 
    process(array_obj_ref_90_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_90_root_address_inst:flowthrough  inputs: " & " read_write_bar_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_buffer) & " array_obj_ref_90_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_90_final_offset) & "outputs: " & " array_obj_ref_90_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_90_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_90_root_address_inst
    process(array_obj_ref_90_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_90_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_90_root_address <= ov(10 downto 0);
      --
    end process;
    -- logger for split-operator ADD_u12_u12_34_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_34_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:ADD_u12_u12_34_inst:started:   inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " addr_buffer = "& Convert_SLV_To_Hex_String(addr_buffer) & " konst_33_wire_constant = "& Convert_SLV_To_Hex_String(konst_33_wire_constant));
          --
        end if; 
        if ADD_u12_u12_34_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:ADD_u12_u12_34_inst:finished:  outputs: " & " addr1_35= "  & Convert_SLV_To_Hex_String(addr1_35));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (0) : ADD_u12_u12_34_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= addr_buffer;
      addr1_35 <= data_out(11 downto 0);
      guard_vector(0)  <= read_write_bar_buffer(0);
      reqL_unguarded(0) <= ADD_u12_u12_34_inst_req_0;
      ADD_u12_u12_34_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_34_inst_req_1;
      ADD_u12_u12_34_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000000000001",
          constant_width => 12,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- logger for split-operator ADD_u12_u12_48_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_48_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:ADD_u12_u12_48_inst:started:   inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " addr_buffer = "& Convert_SLV_To_Hex_String(addr_buffer) & " konst_47_wire_constant = "& Convert_SLV_To_Hex_String(konst_47_wire_constant));
          --
        end if; 
        if ADD_u12_u12_48_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:ADD_u12_u12_48_inst:finished:  outputs: " & " addr2_49= "  & Convert_SLV_To_Hex_String(addr2_49));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (1) : ADD_u12_u12_48_inst 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= addr_buffer;
      addr2_49 <= data_out(11 downto 0);
      guard_vector(0)  <= read_write_bar_buffer(0);
      reqL_unguarded(0) <= ADD_u12_u12_48_inst_req_0;
      ADD_u12_u12_48_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_48_inst_req_1;
      ADD_u12_u12_48_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000000000010",
          constant_width => 12,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- logger for split-operator ADD_u12_u12_62_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_62_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:ADD_u12_u12_62_inst:started:   inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " addr_buffer = "& Convert_SLV_To_Hex_String(addr_buffer) & " konst_61_wire_constant = "& Convert_SLV_To_Hex_String(konst_61_wire_constant));
          --
        end if; 
        if ADD_u12_u12_62_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:ADD_u12_u12_62_inst:finished:  outputs: " & " addr3_63= "  & Convert_SLV_To_Hex_String(addr3_63));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (2) : ADD_u12_u12_62_inst 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= addr_buffer;
      addr3_63 <= data_out(11 downto 0);
      guard_vector(0)  <= read_write_bar_buffer(0);
      reqL_unguarded(0) <= ADD_u12_u12_62_inst_req_0;
      ADD_u12_u12_62_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_62_inst_req_1;
      ADD_u12_u12_62_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_2_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000000000011",
          constant_width => 12,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- logger for split-operator CONCAT_u16_u32_82_inst flow-through 
    process(CONCAT_u16_u32_82_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:CONCAT_u16_u32_82_inst:flowthrough inputs: " & " read_write_bar_63_delayed_6_0_77 (guard)= " & Convert_SLV_To_String(read_write_bar_63_delayed_6_0_77) & " t_read_data3_71 = "& Convert_SLV_To_Hex_String(t_read_data3_71) & " t_read_data2_57 = "& Convert_SLV_To_Hex_String(t_read_data2_57) & " outputs:" & " CONCAT_u16_u32_82_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u16_u32_82_wire));
      --
    end process; 
    -- binary operator CONCAT_u16_u32_82_inst
    process(t_read_data3_71, t_read_data2_57) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(t_read_data3_71, t_read_data2_57, tmp_var);
      CONCAT_u16_u32_82_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u16_u32_85_inst flow-through 
    process(CONCAT_u16_u32_85_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:CONCAT_u16_u32_85_inst:flowthrough inputs: " & " read_write_bar_63_delayed_6_0_77 (guard)= " & Convert_SLV_To_String(read_write_bar_63_delayed_6_0_77) & " t_read_data1_43 = "& Convert_SLV_To_Hex_String(t_read_data1_43) & " t_read_data0_69_delayed_1_0_74 = "& Convert_SLV_To_Hex_String(t_read_data0_69_delayed_1_0_74) & " outputs:" & " CONCAT_u16_u32_85_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u16_u32_85_wire));
      --
    end process; 
    -- binary operator CONCAT_u16_u32_85_inst
    process(t_read_data1_43, t_read_data0_69_delayed_1_0_74) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(t_read_data1_43, t_read_data0_69_delayed_1_0_74, tmp_var);
      CONCAT_u16_u32_85_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u32_u64_86_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if CONCAT_u32_u64_86_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:CONCAT_u32_u64_86_inst:started:   inputs: " & " read_write_bar_63_delayed_6_0_77 (guard)= " & Convert_SLV_To_String(read_write_bar_63_delayed_6_0_77) & " CONCAT_u16_u32_82_wire = "& Convert_SLV_To_Hex_String(CONCAT_u16_u32_82_wire) & " CONCAT_u16_u32_85_wire = "& Convert_SLV_To_Hex_String(CONCAT_u16_u32_85_wire));
          --
        end if; 
        if CONCAT_u32_u64_86_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:CONCAT_u32_u64_86_inst:finished:  outputs: " & " t_read_datal_87= "  & Convert_SLV_To_Hex_String(t_read_datal_87));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (5) : CONCAT_u32_u64_86_inst 
    ApConcat_group_5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_82_wire & CONCAT_u16_u32_85_wire;
      t_read_datal_87 <= data_out(63 downto 0);
      guard_vector(0)  <= read_write_bar_63_delayed_6_0_77(0);
      reqL_unguarded(0) <= CONCAT_u32_u64_86_inst_req_0;
      CONCAT_u32_u64_86_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_86_inst_req_1;
      CONCAT_u32_u64_86_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_5_gI: SplitGuardInterface generic map(name => "ApConcat_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- logger for split-operator array_obj_ref_42_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_42_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_42_load_0:started:   inputs: " & " read_write_bar_36_delayed_1_0_38 (guard)= " & Convert_SLV_To_String(read_write_bar_36_delayed_1_0_38) & " array_obj_ref_42_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_42_word_address_0));
          --
        end if; 
        if array_obj_ref_42_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_42_load_0:finished:  outputs: " & " array_obj_ref_42_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_42_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_28_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_28_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_28_load_0:started:   inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " array_obj_ref_28_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_28_word_address_0));
          --
        end if; 
        if array_obj_ref_28_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_28_load_0:finished:  outputs: " & " array_obj_ref_28_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_28_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_56_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_56_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_56_load_0:started:   inputs: " & " read_write_bar_47_delayed_1_0_52 (guard)= " & Convert_SLV_To_String(read_write_bar_47_delayed_1_0_52) & " array_obj_ref_56_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_56_word_address_0));
          --
        end if; 
        if array_obj_ref_56_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_56_load_0:finished:  outputs: " & " array_obj_ref_56_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_56_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_70_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_70_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_70_load_0:started:   inputs: " & " read_write_bar_58_delayed_1_0_66 (guard)= " & Convert_SLV_To_String(read_write_bar_58_delayed_1_0_66) & " array_obj_ref_70_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_70_word_address_0));
          --
        end if; 
        if array_obj_ref_70_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_70_load_0:finished:  outputs: " & " array_obj_ref_70_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_70_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (0) : array_obj_ref_42_load_0 array_obj_ref_28_load_0 array_obj_ref_56_load_0 array_obj_ref_70_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(43 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => true, 1 => true, 2 => true, 3 => true);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 5, 1 => 5, 2 => 5, 3 => 5);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_42_load_0_req_0,
        array_obj_ref_42_load_0_ack_0,
        array_obj_ref_42_load_0_req_1,
        array_obj_ref_42_load_0_ack_1,
        "array_obj_ref_42_load_0",
        "memory_space_5" ,
        array_obj_ref_42_data_0,
        array_obj_ref_42_word_address_0,
        "array_obj_ref_42_data_0",
        "array_obj_ref_42_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_28_load_0_req_0,
        array_obj_ref_28_load_0_ack_0,
        array_obj_ref_28_load_0_req_1,
        array_obj_ref_28_load_0_ack_1,
        "array_obj_ref_28_load_0",
        "memory_space_5" ,
        array_obj_ref_28_data_0,
        array_obj_ref_28_word_address_0,
        "array_obj_ref_28_data_0",
        "array_obj_ref_28_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_56_load_0_req_0,
        array_obj_ref_56_load_0_ack_0,
        array_obj_ref_56_load_0_req_1,
        array_obj_ref_56_load_0_ack_1,
        "array_obj_ref_56_load_0",
        "memory_space_5" ,
        array_obj_ref_56_data_0,
        array_obj_ref_56_word_address_0,
        "array_obj_ref_56_data_0",
        "array_obj_ref_56_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_70_load_0_req_0,
        array_obj_ref_70_load_0_ack_0,
        array_obj_ref_70_load_0_req_1,
        array_obj_ref_70_load_0_ack_1,
        "array_obj_ref_70_load_0",
        "memory_space_5" ,
        array_obj_ref_70_data_0,
        array_obj_ref_70_word_address_0,
        "array_obj_ref_70_data_0",
        "array_obj_ref_70_word_address_0" -- 
      );
      reqL_unguarded(3) <= array_obj_ref_42_load_0_req_0;
      reqL_unguarded(2) <= array_obj_ref_28_load_0_req_0;
      reqL_unguarded(1) <= array_obj_ref_56_load_0_req_0;
      reqL_unguarded(0) <= array_obj_ref_70_load_0_req_0;
      array_obj_ref_42_load_0_ack_0 <= ackL_unguarded(3);
      array_obj_ref_28_load_0_ack_0 <= ackL_unguarded(2);
      array_obj_ref_56_load_0_ack_0 <= ackL_unguarded(1);
      array_obj_ref_70_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= array_obj_ref_42_load_0_req_1;
      reqR_unguarded(2) <= array_obj_ref_28_load_0_req_1;
      reqR_unguarded(1) <= array_obj_ref_56_load_0_req_1;
      reqR_unguarded(0) <= array_obj_ref_70_load_0_req_1;
      array_obj_ref_42_load_0_ack_1 <= ackR_unguarded(3);
      array_obj_ref_28_load_0_ack_1 <= ackR_unguarded(2);
      array_obj_ref_56_load_0_ack_1 <= ackR_unguarded(1);
      array_obj_ref_70_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_write_bar_58_delayed_1_0_66(0);
      guard_vector(1)  <= read_write_bar_47_delayed_1_0_52(0);
      guard_vector(2)  <= read_write_bar_buffer(0);
      guard_vector(3)  <= read_write_bar_36_delayed_1_0_38(0);
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_42_word_address_0 & array_obj_ref_28_word_address_0 & array_obj_ref_56_word_address_0 & array_obj_ref_70_word_address_0;
      array_obj_ref_42_data_0 <= data_out(63 downto 48);
      array_obj_ref_28_data_0 <= data_out(47 downto 32);
      array_obj_ref_56_data_0 <= data_out(31 downto 16);
      array_obj_ref_70_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 11,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(10 downto 0),
          mtag => memory_space_5_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(15 downto 0),
          mtag => memory_space_5_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logger for split-operator array_obj_ref_90_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_90_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_90_store_0:started:   inputs: " & " read_write_bar_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_buffer) & " array_obj_ref_90_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_90_word_address_0) & " array_obj_ref_90_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_90_data_0));
          --
        end if; 
        if array_obj_ref_90_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_90_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_90_store_0_req_0,
      array_obj_ref_90_store_0_ack_0,
      array_obj_ref_90_store_0_req_1,
      array_obj_ref_90_store_0_ack_1,
      "array_obj_ref_90_store_0",
      "memory_space_5" ,
      array_obj_ref_90_data_0,
      array_obj_ref_90_word_address_0,
      "array_obj_ref_90_data_0",
      "array_obj_ref_90_word_address_0" -- 
    );
    -- shared store operator group (0) : array_obj_ref_90_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_90_store_0_req_0;
      array_obj_ref_90_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_90_store_0_req_1;
      array_obj_ref_90_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_write_bar_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_90_word_address_0;
      data_in <= array_obj_ref_90_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 11,
        data_width => 16,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(10 downto 0),
          mdata => memory_space_5_sr_data(15 downto 0),
          mtag => memory_space_5_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end accessMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity accessMem_v is -- 
  generic (tag_length : integer); 
  port ( -- 
    read_write_bar : in  std_logic_vector(0 downto 0);
    addr : in  std_logic_vector(11 downto 0);
    write_data : in  std_logic_vector(15 downto 0);
    read_datal : out  std_logic_vector(63 downto 0);
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(10 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessMem_v;
architecture accessMem_v_arch of accessMem_v is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 29)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal read_write_bar_buffer :  std_logic_vector(0 downto 0);
  signal read_write_bar_update_enable: Boolean;
  signal addr_buffer :  std_logic_vector(11 downto 0);
  signal addr_update_enable: Boolean;
  signal write_data_buffer :  std_logic_vector(15 downto 0);
  signal write_data_update_enable: Boolean;
  -- output port buffer signals
  signal read_datal_buffer :  std_logic_vector(63 downto 0);
  signal read_datal_update_enable: Boolean;
  signal accessMem_v_CP_553_start: Boolean;
  signal accessMem_v_CP_553_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ADD_u12_u12_157_inst_ack_1 : boolean;
  signal ADD_u12_u12_157_inst_req_1 : boolean;
  signal ADD_u12_u12_157_inst_ack_0 : boolean;
  signal ADD_u12_u12_157_inst_req_0 : boolean;
  signal array_obj_ref_151_load_0_ack_1 : boolean;
  signal array_obj_ref_151_load_0_req_1 : boolean;
  signal array_obj_ref_151_load_0_ack_0 : boolean;
  signal array_obj_ref_151_load_0_req_0 : boolean;
  signal array_obj_ref_165_load_0_ack_1 : boolean;
  signal array_obj_ref_165_load_0_req_1 : boolean;
  signal W_read_write_bar_146_delayed_1_0_159_inst_ack_1 : boolean;
  signal W_read_write_bar_168_delayed_1_0_187_inst_ack_1 : boolean;
  signal array_obj_ref_165_load_0_ack_0 : boolean;
  signal array_obj_ref_165_load_0_req_0 : boolean;
  signal W_read_write_bar_168_delayed_1_0_187_inst_req_1 : boolean;
  signal W_read_write_bar_146_delayed_1_0_159_inst_req_1 : boolean;
  signal ADD_u12_u12_185_inst_ack_1 : boolean;
  signal W_read_write_bar_157_delayed_1_0_173_inst_ack_1 : boolean;
  signal ADD_u12_u12_185_inst_req_1 : boolean;
  signal W_read_write_bar_157_delayed_1_0_173_inst_req_1 : boolean;
  signal W_read_write_bar_168_delayed_1_0_187_inst_req_0 : boolean;
  signal W_read_write_bar_168_delayed_1_0_187_inst_ack_0 : boolean;
  signal ADD_u12_u12_185_inst_req_0 : boolean;
  signal ADD_u12_u12_185_inst_ack_0 : boolean;
  signal W_read_write_bar_157_delayed_1_0_173_inst_ack_0 : boolean;
  signal W_read_write_bar_157_delayed_1_0_173_inst_req_0 : boolean;
  signal ADD_u12_u12_171_inst_ack_0 : boolean;
  signal ADD_u12_u12_171_inst_req_0 : boolean;
  signal W_read_write_bar_146_delayed_1_0_159_inst_ack_0 : boolean;
  signal W_read_write_bar_146_delayed_1_0_159_inst_req_0 : boolean;
  signal array_obj_ref_179_load_0_ack_1 : boolean;
  signal array_obj_ref_179_load_0_req_1 : boolean;
  signal ADD_u12_u12_171_inst_ack_1 : boolean;
  signal ADD_u12_u12_171_inst_req_1 : boolean;
  signal array_obj_ref_179_load_0_ack_0 : boolean;
  signal array_obj_ref_179_load_0_req_0 : boolean;
  signal array_obj_ref_193_load_0_req_0 : boolean;
  signal array_obj_ref_193_load_0_ack_0 : boolean;
  signal array_obj_ref_193_load_0_req_1 : boolean;
  signal array_obj_ref_193_load_0_ack_1 : boolean;
  signal W_read_write_bar_173_delayed_6_0_195_inst_req_0 : boolean;
  signal W_read_write_bar_173_delayed_6_0_195_inst_ack_0 : boolean;
  signal W_read_write_bar_173_delayed_6_0_195_inst_req_1 : boolean;
  signal W_read_write_bar_173_delayed_6_0_195_inst_ack_1 : boolean;
  signal W_t_read_data0_179_delayed_1_0_198_inst_req_0 : boolean;
  signal W_t_read_data0_179_delayed_1_0_198_inst_ack_0 : boolean;
  signal W_t_read_data0_179_delayed_1_0_198_inst_req_1 : boolean;
  signal W_t_read_data0_179_delayed_1_0_198_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_209_inst_req_0 : boolean;
  signal CONCAT_u32_u64_209_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_209_inst_req_1 : boolean;
  signal CONCAT_u32_u64_209_inst_ack_1 : boolean;
  signal array_obj_ref_213_store_0_req_0 : boolean;
  signal array_obj_ref_213_store_0_ack_0 : boolean;
  signal array_obj_ref_213_store_0_req_1 : boolean;
  signal array_obj_ref_213_store_0_ack_1 : boolean;
  signal W_read_write_bar_189_delayed_7_0_216_inst_req_0 : boolean;
  signal W_read_write_bar_189_delayed_7_0_216_inst_ack_0 : boolean;
  signal W_read_write_bar_189_delayed_7_0_216_inst_req_1 : boolean;
  signal W_read_write_bar_189_delayed_7_0_216_inst_ack_1 : boolean;
  signal MUX_223_inst_req_0 : boolean;
  signal MUX_223_inst_ack_0 : boolean;
  signal MUX_223_inst_req_1 : boolean;
  signal MUX_223_inst_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessMem_v_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 29) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= read_write_bar;
  read_write_bar_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(12 downto 1) <= addr;
  addr_buffer <= in_buffer_data_out(12 downto 1);
  in_buffer_data_in(28 downto 13) <= write_data;
  write_data_buffer <= in_buffer_data_out(28 downto 13);
  in_buffer_data_in(tag_length + 28 downto 29) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 28 downto 29);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 4) := (0 => 14,1 => 14,2 => 14,3 => 1,4 => 14);
    constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 14);
    constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 5); -- 
  begin -- 
    preds <= read_write_bar_update_enable & addr_update_enable & write_data_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessMem_v_CP_553_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessMem_v_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= read_datal_buffer;
  read_datal <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 14,1 => 1,2 => 14);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMem_v_CP_553_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  read_datal_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 29) := "read_datal_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_read_datal_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => read_datal_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 14,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 14,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessMem_v_CP_553_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 14,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMem_v_CP_553_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,accessMem_v_CP_553_start,"accessMem_v cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,accessMem_v_CP_553_symbol, "accessMem_v cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessMem_v_CP_553: Block -- control-path 
    signal accessMem_v_CP_553_elements: BooleanArray(79 downto 0);
    -- 
  begin -- 
    accessMem_v_CP_553_elements(0) <= accessMem_v_CP_553_start;
    accessMem_v_CP_553_symbol <= accessMem_v_CP_553_elements(79);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	6 
    -- CP-element group 1: 	10 
    -- CP-element group 1: 	14 
    -- CP-element group 1: 	22 
    -- CP-element group 1: 	26 
    -- CP-element group 1: 	34 
    -- CP-element group 1: 	38 
    -- CP-element group 1: 	46 
    -- CP-element group 1: 	58 
    -- CP-element group 1: 	62 
    -- CP-element group 1:  members (53) 
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_index_scale_0/$exit
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_index_scale_0/$entry
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_index_resize_0/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_word_addrgen/root_register_ack
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_word_addrgen/root_register_req
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_word_addrgen/$exit
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_word_addrgen/$entry
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_base_plus_offset/sum_rename_ack
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_base_plus_offset/sum_rename_req
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_base_plus_offset/$exit
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_base_plus_offset/$entry
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_final_index_sum_regn/ack
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_final_index_sum_regn/req
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_final_index_sum_regn/$exit
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_final_index_sum_regn/$entry
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_index_scale_0/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_index_scale_0/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_index_resize_0/index_resize_req
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_index_resize_0/$exit
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_index_resize_0/$entry
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_index_computed_0
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_index_scaled_0
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_index_resized_0
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_offset_calculated
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_root_address_calculated
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_word_address_calculated
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/$entry
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_word_address_calculated
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_root_address_calculated
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_offset_calculated
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_index_resized_0
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_index_scaled_0
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_index_computed_0
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_index_resize_0/$entry
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_index_resize_0/$exit
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_index_resize_0/index_resize_req
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_index_resize_0/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_index_scale_0/$entry
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_index_scale_0/$exit
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_index_scale_0/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_index_scale_0/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_final_index_sum_regn/$entry
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_final_index_sum_regn/$exit
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_final_index_sum_regn/req
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_final_index_sum_regn/ack
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_base_plus_offset/$entry
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_base_plus_offset/$exit
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_base_plus_offset/sum_rename_req
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_base_plus_offset/sum_rename_ack
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_word_addrgen/$entry
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_word_addrgen/$exit
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_word_addrgen/root_register_req
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_v_CP_553_elements(1) <= accessMem_v_CP_553_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	36 
    -- CP-element group 2: 	40 
    -- CP-element group 2: 	48 
    -- CP-element group 2: 	60 
    -- CP-element group 2: 	64 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	75 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_152_to_assign_stmt_224/read_write_bar_update_enable_out
      -- CP-element group 2: 	 assign_stmt_152_to_assign_stmt_224/read_write_bar_update_enable
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_v_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 30) := "accessMem_v_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(8) & accessMem_v_CP_553_elements(12) & accessMem_v_CP_553_elements(16) & accessMem_v_CP_553_elements(24) & accessMem_v_CP_553_elements(28) & accessMem_v_CP_553_elements(36) & accessMem_v_CP_553_elements(40) & accessMem_v_CP_553_elements(48) & accessMem_v_CP_553_elements(60) & accessMem_v_CP_553_elements(64);
      gj_accessMem_v_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	8 
    -- CP-element group 3: 	12 
    -- CP-element group 3: 	24 
    -- CP-element group 3: 	36 
    -- CP-element group 3: 	60 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	76 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_152_to_assign_stmt_224/addr_update_enable_out
      -- CP-element group 3: 	 assign_stmt_152_to_assign_stmt_224/addr_update_enable
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_v_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "accessMem_v_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(8) & accessMem_v_CP_553_elements(12) & accessMem_v_CP_553_elements(24) & accessMem_v_CP_553_elements(36) & accessMem_v_CP_553_elements(60);
      gj_accessMem_v_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	60 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	77 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_152_to_assign_stmt_224/write_data_update_enable_out
      -- CP-element group 4: 	 assign_stmt_152_to_assign_stmt_224/write_data_update_enable
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_v_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "accessMem_v_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMem_v_CP_553_elements(60);
      gj_accessMem_v_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	78 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	67 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_152_to_assign_stmt_224/read_datal_update_enable_in
      -- CP-element group 5: 	 assign_stmt_152_to_assign_stmt_224/read_datal_update_enable
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_v_CP_553_elements(5) <= accessMem_v_CP_553_elements(78);
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	1 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	8 
    -- CP-element group 6: 	60 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (5) 
      -- CP-element group 6: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_Sample/word_access_start/word_0/rr
      -- CP-element group 6: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_Sample/word_access_start/word_0/$entry
      -- CP-element group 6: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_Sample/word_access_start/$entry
      -- CP-element group 6: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_Sample/$entry
      -- CP-element group 6: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_sample_start_
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:array_obj_ref_151_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(6), ack => array_obj_ref_151_load_0_req_0); -- 
    accessMem_v_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 14,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 30) := "accessMem_v_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(1) & accessMem_v_CP_553_elements(8) & accessMem_v_CP_553_elements(60);
      gj_accessMem_v_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: marked-predecessors 
    -- CP-element group 7: 	9 
    -- CP-element group 7: 	52 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	9 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_Update/word_access_complete/word_0/cr
      -- CP-element group 7: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_Update/word_access_complete/word_0/$entry
      -- CP-element group 7: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_Update/word_access_complete/$entry
      -- CP-element group 7: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_Update/$entry
      -- CP-element group 7: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_update_start_
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:array_obj_ref_151_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(7), ack => array_obj_ref_151_load_0_req_1); -- 
    accessMem_v_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "accessMem_v_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(9) & accessMem_v_CP_553_elements(52);
      gj_accessMem_v_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	70 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: 	3 
    -- CP-element group 8: 	6 
    -- CP-element group 8:  members (5) 
      -- CP-element group 8: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_Sample/word_access_start/word_0/ra
      -- CP-element group 8: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_Sample/word_access_start/word_0/$exit
      -- CP-element group 8: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_Sample/word_access_start/$exit
      -- CP-element group 8: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_Sample/$exit
      -- CP-element group 8: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_sample_completed_
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:array_obj_ref_151_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_151_load_0_ack_0, ack => accessMem_v_CP_553_elements(8)); -- 
    -- CP-element group 9:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	7 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	50 
    -- CP-element group 9: marked-successors 
    -- CP-element group 9: 	7 
    -- CP-element group 9:  members (9) 
      -- CP-element group 9: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_Update/array_obj_ref_151_Merge/$exit
      -- CP-element group 9: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_Update/array_obj_ref_151_Merge/merge_ack
      -- CP-element group 9: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_Update/array_obj_ref_151_Merge/merge_req
      -- CP-element group 9: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_Update/array_obj_ref_151_Merge/$entry
      -- CP-element group 9: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_Update/word_access_complete/word_0/ca
      -- CP-element group 9: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_Update/word_access_complete/word_0/$exit
      -- CP-element group 9: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_Update/word_access_complete/$exit
      -- CP-element group 9: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_Update/$exit
      -- CP-element group 9: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_update_completed_
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(9) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:array_obj_ref_151_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_151_load_0_ack_1, ack => accessMem_v_CP_553_elements(9)); -- 
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	1 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_157_Sample/rr
      -- CP-element group 10: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_157_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_157_sample_start_
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:ADD_u12_u12_157_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(10), ack => ADD_u12_u12_157_inst_req_0); -- 
    accessMem_v_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 14,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(1) & accessMem_v_CP_553_elements(12);
      gj_accessMem_v_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	13 
    -- CP-element group 11: 	20 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_157_Update/cr
      -- CP-element group 11: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_157_Update/$entry
      -- CP-element group 11: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_157_update_start_
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:ADD_u12_u12_157_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(11), ack => ADD_u12_u12_157_inst_req_1); -- 
    accessMem_v_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(13) & accessMem_v_CP_553_elements(20);
      gj_accessMem_v_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: 	3 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_157_Sample/ra
      -- CP-element group 12: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_157_Sample/$exit
      -- CP-element group 12: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_157_sample_completed_
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:ADD_u12_u12_157_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_157_inst_ack_0, ack => accessMem_v_CP_553_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	18 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	11 
    -- CP-element group 13:  members (29) 
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_final_index_sum_regn/ack
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_157_Update/ca
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_157_Update/$exit
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_157_update_completed_
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_final_index_sum_regn/req
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_index_resize_0/$entry
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_index_scale_0/$exit
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_root_address_calculated
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_final_index_sum_regn/$exit
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_word_address_calculated
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_final_index_sum_regn/$entry
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_index_scale_0/scale_rename_ack
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_index_scale_0/scale_rename_req
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_index_computed_0
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_index_scale_0/$entry
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_word_addrgen/root_register_ack
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_word_addrgen/root_register_req
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_word_addrgen/$exit
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_word_addrgen/$entry
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_index_scaled_0
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_index_resize_0/index_resize_ack
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_base_plus_offset/sum_rename_ack
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_base_plus_offset/sum_rename_req
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_base_plus_offset/$exit
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_index_resize_0/index_resize_req
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_base_plus_offset/$entry
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_index_resized_0
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_offset_calculated
      -- CP-element group 13: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_index_resize_0/$exit
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:ADD_u12_u12_157_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_157_inst_ack_1, ack => accessMem_v_CP_553_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	1 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_161_sample_start_
      -- CP-element group 14: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_161_Sample/$entry
      -- CP-element group 14: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_161_Sample/req
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_read_write_bar_146_delayed_1_0_159_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(14), ack => W_read_write_bar_146_delayed_1_0_159_inst_req_0); -- 
    accessMem_v_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 14,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(1) & accessMem_v_CP_553_elements(16);
      gj_accessMem_v_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	20 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_161_update_start_
      -- CP-element group 15: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_161_Update/req
      -- CP-element group 15: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_161_Update/$entry
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_read_write_bar_146_delayed_1_0_159_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(15), ack => W_read_write_bar_146_delayed_1_0_159_inst_req_1); -- 
    accessMem_v_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(17) & accessMem_v_CP_553_elements(20);
      gj_accessMem_v_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_161_sample_completed_
      -- CP-element group 16: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_161_Sample/$exit
      -- CP-element group 16: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_161_Sample/ack
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_read_write_bar_146_delayed_1_0_159_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_146_delayed_1_0_159_inst_ack_0, ack => accessMem_v_CP_553_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	15 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_161_update_completed_
      -- CP-element group 17: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_161_Update/ack
      -- CP-element group 17: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_161_Update/$exit
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_read_write_bar_146_delayed_1_0_159_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_146_delayed_1_0_159_inst_ack_1, ack => accessMem_v_CP_553_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	13 
    -- CP-element group 18: 	17 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: 	60 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (5) 
      -- CP-element group 18: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_sample_start_
      -- CP-element group 18: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_Sample/word_access_start/$entry
      -- CP-element group 18: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_Sample/word_access_start/word_0/rr
      -- CP-element group 18: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_Sample/word_access_start/word_0/$entry
      -- CP-element group 18: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_Sample/$entry
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:array_obj_ref_165_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(18), ack => array_obj_ref_165_load_0_req_0); -- 
    accessMem_v_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(13) & accessMem_v_CP_553_elements(17) & accessMem_v_CP_553_elements(20) & accessMem_v_CP_553_elements(60);
      gj_accessMem_v_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	21 
    -- CP-element group 19: 	56 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_Update/word_access_complete/word_0/cr
      -- CP-element group 19: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_Update/word_access_complete/word_0/$entry
      -- CP-element group 19: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_Update/word_access_complete/$entry
      -- CP-element group 19: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_Update/$entry
      -- CP-element group 19: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_update_start_
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:array_obj_ref_165_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(19), ack => array_obj_ref_165_load_0_req_1); -- 
    accessMem_v_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(21) & accessMem_v_CP_553_elements(56);
      gj_accessMem_v_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	71 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	11 
    -- CP-element group 20: 	15 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (5) 
      -- CP-element group 20: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_Sample/$exit
      -- CP-element group 20: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_Sample/word_access_start/word_0/ra
      -- CP-element group 20: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_Sample/word_access_start/word_0/$exit
      -- CP-element group 20: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_Sample/word_access_start/$exit
      -- CP-element group 20: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_sample_completed_
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:array_obj_ref_165_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_165_load_0_ack_0, ack => accessMem_v_CP_553_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	54 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	19 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_Update/array_obj_ref_165_Merge/merge_ack
      -- CP-element group 21: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_Update/array_obj_ref_165_Merge/merge_req
      -- CP-element group 21: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_Update/array_obj_ref_165_Merge/$exit
      -- CP-element group 21: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_Update/array_obj_ref_165_Merge/$entry
      -- CP-element group 21: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_Update/word_access_complete/word_0/ca
      -- CP-element group 21: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_Update/word_access_complete/word_0/$exit
      -- CP-element group 21: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_Update/word_access_complete/$exit
      -- CP-element group 21: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_Update/$exit
      -- CP-element group 21: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_update_completed_
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:array_obj_ref_165_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_165_load_0_ack_1, ack => accessMem_v_CP_553_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	1 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	24 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_171_Sample/$entry
      -- CP-element group 22: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_171_sample_start_
      -- CP-element group 22: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_171_Sample/rr
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:ADD_u12_u12_171_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(22), ack => ADD_u12_u12_171_inst_req_0); -- 
    accessMem_v_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 14,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(1) & accessMem_v_CP_553_elements(24);
      gj_accessMem_v_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: 	32 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_171_update_start_
      -- CP-element group 23: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_171_Update/$entry
      -- CP-element group 23: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_171_Update/cr
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:ADD_u12_u12_171_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(23), ack => ADD_u12_u12_171_inst_req_1); -- 
    accessMem_v_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(25) & accessMem_v_CP_553_elements(32);
      gj_accessMem_v_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: 	3 
    -- CP-element group 24: 	22 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_171_Sample/$exit
      -- CP-element group 24: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_171_sample_completed_
      -- CP-element group 24: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_171_Sample/ra
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:ADD_u12_u12_171_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_171_inst_ack_0, ack => accessMem_v_CP_553_elements(24)); -- 
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	30 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	23 
    -- CP-element group 25:  members (29) 
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_index_resize_0/$entry
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_index_resize_0/$exit
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_index_resized_0
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_index_computed_0
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_offset_calculated
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_index_scaled_0
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_root_address_calculated
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_word_address_calculated
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_171_update_completed_
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_171_Update/$exit
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_word_addrgen/root_register_ack
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_word_addrgen/root_register_req
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_word_addrgen/$exit
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_word_addrgen/$entry
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_base_plus_offset/sum_rename_ack
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_base_plus_offset/sum_rename_req
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_base_plus_offset/$entry
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_base_plus_offset/$exit
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_final_index_sum_regn/ack
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_final_index_sum_regn/req
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_final_index_sum_regn/$entry
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_final_index_sum_regn/$exit
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_171_Update/ca
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_index_scale_0/scale_rename_ack
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_index_scale_0/scale_rename_req
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_index_scale_0/$entry
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_index_scale_0/$exit
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_index_resize_0/index_resize_ack
      -- CP-element group 25: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_index_resize_0/index_resize_req
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:ADD_u12_u12_171_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_171_inst_ack_1, ack => accessMem_v_CP_553_elements(25)); -- 
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	1 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	28 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_175_sample_start_
      -- CP-element group 26: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_175_Sample/$entry
      -- CP-element group 26: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_175_Sample/req
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_read_write_bar_157_delayed_1_0_173_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(26), ack => W_read_write_bar_157_delayed_1_0_173_inst_req_0); -- 
    accessMem_v_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 14,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(1) & accessMem_v_CP_553_elements(28);
      gj_accessMem_v_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: 	32 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_175_update_start_
      -- CP-element group 27: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_175_Update/req
      -- CP-element group 27: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_175_Update/$entry
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_read_write_bar_157_delayed_1_0_173_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(27), ack => W_read_write_bar_157_delayed_1_0_173_inst_req_1); -- 
    accessMem_v_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(29) & accessMem_v_CP_553_elements(32);
      gj_accessMem_v_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: 	26 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_175_sample_completed_
      -- CP-element group 28: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_175_Sample/$exit
      -- CP-element group 28: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_175_Sample/ack
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_read_write_bar_157_delayed_1_0_173_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_157_delayed_1_0_173_inst_ack_0, ack => accessMem_v_CP_553_elements(28)); -- 
    -- CP-element group 29:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_175_update_completed_
      -- CP-element group 29: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_175_Update/ack
      -- CP-element group 29: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_175_Update/$exit
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_read_write_bar_157_delayed_1_0_173_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_157_delayed_1_0_173_inst_ack_1, ack => accessMem_v_CP_553_elements(29)); -- 
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	25 
    -- CP-element group 30: 	29 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: 	60 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (5) 
      -- CP-element group 30: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_sample_start_
      -- CP-element group 30: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_Sample/word_access_start/word_0/$entry
      -- CP-element group 30: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_Sample/word_access_start/$entry
      -- CP-element group 30: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_Sample/$entry
      -- CP-element group 30: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:array_obj_ref_179_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(30), ack => array_obj_ref_179_load_0_req_0); -- 
    accessMem_v_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(25) & accessMem_v_CP_553_elements(29) & accessMem_v_CP_553_elements(32) & accessMem_v_CP_553_elements(60);
      gj_accessMem_v_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: 	56 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (5) 
      -- CP-element group 31: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_update_start_
      -- CP-element group 31: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_Update/word_access_complete/word_0/cr
      -- CP-element group 31: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_Update/word_access_complete/word_0/$entry
      -- CP-element group 31: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_Update/word_access_complete/$entry
      -- CP-element group 31: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_Update/$entry
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:array_obj_ref_179_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(31), ack => array_obj_ref_179_load_0_req_1); -- 
    accessMem_v_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(33) & accessMem_v_CP_553_elements(56);
      gj_accessMem_v_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	72 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	23 
    -- CP-element group 32: 	27 
    -- CP-element group 32: 	30 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_sample_completed_
      -- CP-element group 32: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_Sample/word_access_start/word_0/$exit
      -- CP-element group 32: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_Sample/word_access_start/$exit
      -- CP-element group 32: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_Sample/$exit
      -- CP-element group 32: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:array_obj_ref_179_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_179_load_0_ack_0, ack => accessMem_v_CP_553_elements(32)); -- 
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	54 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (9) 
      -- CP-element group 33: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_update_completed_
      -- CP-element group 33: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_Update/array_obj_ref_179_Merge/merge_ack
      -- CP-element group 33: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_Update/array_obj_ref_179_Merge/merge_req
      -- CP-element group 33: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_Update/array_obj_ref_179_Merge/$exit
      -- CP-element group 33: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_Update/array_obj_ref_179_Merge/$entry
      -- CP-element group 33: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_Update/word_access_complete/word_0/ca
      -- CP-element group 33: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_Update/word_access_complete/word_0/$exit
      -- CP-element group 33: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_Update/$exit
      -- CP-element group 33: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_Update/word_access_complete/$exit
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:array_obj_ref_179_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_179_load_0_ack_1, ack => accessMem_v_CP_553_elements(33)); -- 
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	1 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_185_sample_start_
      -- CP-element group 34: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_185_Sample/$entry
      -- CP-element group 34: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_185_Sample/rr
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:ADD_u12_u12_185_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(34), ack => ADD_u12_u12_185_inst_req_0); -- 
    accessMem_v_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 14,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(1) & accessMem_v_CP_553_elements(36);
      gj_accessMem_v_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	37 
    -- CP-element group 35: 	44 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_185_update_start_
      -- CP-element group 35: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_185_Update/cr
      -- CP-element group 35: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_185_Update/$entry
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:ADD_u12_u12_185_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(35), ack => ADD_u12_u12_185_inst_req_1); -- 
    accessMem_v_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(37) & accessMem_v_CP_553_elements(44);
      gj_accessMem_v_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	2 
    -- CP-element group 36: 	3 
    -- CP-element group 36: 	34 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_185_sample_completed_
      -- CP-element group 36: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_185_Sample/ra
      -- CP-element group 36: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_185_Sample/$exit
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(36) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:ADD_u12_u12_185_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_185_inst_ack_0, ack => accessMem_v_CP_553_elements(36)); -- 
    -- CP-element group 37:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	42 
    -- CP-element group 37: marked-successors 
    -- CP-element group 37: 	35 
    -- CP-element group 37:  members (29) 
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_index_resize_0/$entry
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_index_resize_0/$exit
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_word_address_calculated
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_root_address_calculated
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_index_resized_0
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_index_scaled_0
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_offset_calculated
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_index_resize_0/index_resize_req
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_index_resize_0/index_resize_ack
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_index_computed_0
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_index_scale_0/$entry
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_index_scale_0/$exit
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_185_Update/ca
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_185_Update/$exit
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/ADD_u12_u12_185_update_completed_
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_index_scale_0/scale_rename_req
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_index_scale_0/scale_rename_ack
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_final_index_sum_regn/$entry
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_final_index_sum_regn/$exit
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_final_index_sum_regn/req
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_final_index_sum_regn/ack
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_base_plus_offset/$entry
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_base_plus_offset/$exit
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_base_plus_offset/sum_rename_req
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_base_plus_offset/sum_rename_ack
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_word_addrgen/$entry
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_word_addrgen/$exit
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_word_addrgen/root_register_req
      -- CP-element group 37: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:ADD_u12_u12_185_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_185_inst_ack_1, ack => accessMem_v_CP_553_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	1 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	40 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_189_sample_start_
      -- CP-element group 38: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_189_Sample/req
      -- CP-element group 38: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_189_Sample/$entry
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(38) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_read_write_bar_168_delayed_1_0_187_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(38), ack => W_read_write_bar_168_delayed_1_0_187_inst_req_0); -- 
    accessMem_v_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 14,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(1) & accessMem_v_CP_553_elements(40);
      gj_accessMem_v_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: 	44 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_189_update_start_
      -- CP-element group 39: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_189_Update/req
      -- CP-element group 39: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_189_Update/$entry
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_read_write_bar_168_delayed_1_0_187_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(39), ack => W_read_write_bar_168_delayed_1_0_187_inst_req_1); -- 
    accessMem_v_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(41) & accessMem_v_CP_553_elements(44);
      gj_accessMem_v_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	2 
    -- CP-element group 40: 	38 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_189_Sample/ack
      -- CP-element group 40: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_189_Sample/$exit
      -- CP-element group 40: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_189_sample_completed_
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(40) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_read_write_bar_168_delayed_1_0_187_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_168_delayed_1_0_187_inst_ack_0, ack => accessMem_v_CP_553_elements(40)); -- 
    -- CP-element group 41:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	39 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_189_update_completed_
      -- CP-element group 41: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_189_Update/ack
      -- CP-element group 41: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_189_Update/$exit
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(41) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_read_write_bar_168_delayed_1_0_187_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_168_delayed_1_0_187_inst_ack_1, ack => accessMem_v_CP_553_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	37 
    -- CP-element group 42: 	41 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: 	60 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_sample_start_
      -- CP-element group 42: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_Sample/$entry
      -- CP-element group 42: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_Sample/word_access_start/$entry
      -- CP-element group 42: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_Sample/word_access_start/word_0/$entry
      -- CP-element group 42: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(42) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:array_obj_ref_193_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(42), ack => array_obj_ref_193_load_0_req_0); -- 
    accessMem_v_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(37) & accessMem_v_CP_553_elements(41) & accessMem_v_CP_553_elements(44) & accessMem_v_CP_553_elements(60);
      gj_accessMem_v_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	45 
    -- CP-element group 43: 	56 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (5) 
      -- CP-element group 43: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_update_start_
      -- CP-element group 43: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_Update/$entry
      -- CP-element group 43: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_Update/word_access_complete/$entry
      -- CP-element group 43: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_Update/word_access_complete/word_0/$entry
      -- CP-element group 43: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(43) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:array_obj_ref_193_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(43), ack => array_obj_ref_193_load_0_req_1); -- 
    accessMem_v_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(45) & accessMem_v_CP_553_elements(56);
      gj_accessMem_v_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	73 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	35 
    -- CP-element group 44: 	39 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (5) 
      -- CP-element group 44: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_sample_completed_
      -- CP-element group 44: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_Sample/$exit
      -- CP-element group 44: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_Sample/word_access_start/$exit
      -- CP-element group 44: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_Sample/word_access_start/word_0/$exit
      -- CP-element group 44: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(44) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:array_obj_ref_193_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_193_load_0_ack_0, ack => accessMem_v_CP_553_elements(44)); -- 
    -- CP-element group 45:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	54 
    -- CP-element group 45: marked-successors 
    -- CP-element group 45: 	43 
    -- CP-element group 45:  members (9) 
      -- CP-element group 45: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_update_completed_
      -- CP-element group 45: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_Update/$exit
      -- CP-element group 45: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_Update/word_access_complete/$exit
      -- CP-element group 45: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_Update/word_access_complete/word_0/$exit
      -- CP-element group 45: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_Update/word_access_complete/word_0/ca
      -- CP-element group 45: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_Update/array_obj_ref_193_Merge/$entry
      -- CP-element group 45: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_Update/array_obj_ref_193_Merge/$exit
      -- CP-element group 45: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_Update/array_obj_ref_193_Merge/merge_req
      -- CP-element group 45: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_Update/array_obj_ref_193_Merge/merge_ack
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(45) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:array_obj_ref_193_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_193_load_0_ack_1, ack => accessMem_v_CP_553_elements(45)); -- 
    -- CP-element group 46:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	1 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	48 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_197_sample_start_
      -- CP-element group 46: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_197_Sample/$entry
      -- CP-element group 46: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_197_Sample/req
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(46) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_read_write_bar_173_delayed_6_0_195_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(46), ack => W_read_write_bar_173_delayed_6_0_195_inst_req_0); -- 
    accessMem_v_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 14,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(1) & accessMem_v_CP_553_elements(48);
      gj_accessMem_v_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	49 
    -- CP-element group 47: 	56 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_197_update_start_
      -- CP-element group 47: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_197_Update/$entry
      -- CP-element group 47: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_197_Update/req
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(47) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_read_write_bar_173_delayed_6_0_195_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(47), ack => W_read_write_bar_173_delayed_6_0_195_inst_req_1); -- 
    accessMem_v_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(49) & accessMem_v_CP_553_elements(56);
      gj_accessMem_v_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: marked-successors 
    -- CP-element group 48: 	2 
    -- CP-element group 48: 	46 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_197_sample_completed_
      -- CP-element group 48: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_197_Sample/$exit
      -- CP-element group 48: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_197_Sample/ack
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(48) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_read_write_bar_173_delayed_6_0_195_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_173_delayed_6_0_195_inst_ack_0, ack => accessMem_v_CP_553_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	54 
    -- CP-element group 49: marked-successors 
    -- CP-element group 49: 	47 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_197_update_completed_
      -- CP-element group 49: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_197_Update/$exit
      -- CP-element group 49: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_197_Update/ack
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(49) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_read_write_bar_173_delayed_6_0_195_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_173_delayed_6_0_195_inst_ack_1, ack => accessMem_v_CP_553_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	9 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	52 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_200_sample_start_
      -- CP-element group 50: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_200_Sample/$entry
      -- CP-element group 50: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_200_Sample/req
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(50) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_t_read_data0_179_delayed_1_0_198_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(50), ack => W_t_read_data0_179_delayed_1_0_198_inst_req_0); -- 
    accessMem_v_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(9) & accessMem_v_CP_553_elements(52);
      gj_accessMem_v_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	53 
    -- CP-element group 51: 	56 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_200_update_start_
      -- CP-element group 51: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_200_Update/$entry
      -- CP-element group 51: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_200_Update/req
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(51) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_t_read_data0_179_delayed_1_0_198_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(51), ack => W_t_read_data0_179_delayed_1_0_198_inst_req_1); -- 
    accessMem_v_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(53) & accessMem_v_CP_553_elements(56);
      gj_accessMem_v_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	7 
    -- CP-element group 52: 	50 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_200_sample_completed_
      -- CP-element group 52: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_200_Sample/$exit
      -- CP-element group 52: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_200_Sample/ack
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(52) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_t_read_data0_179_delayed_1_0_198_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_t_read_data0_179_delayed_1_0_198_inst_ack_0, ack => accessMem_v_CP_553_elements(52)); -- 
    -- CP-element group 53:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53: marked-successors 
    -- CP-element group 53: 	51 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_200_update_completed_
      -- CP-element group 53: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_200_Update/$exit
      -- CP-element group 53: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_200_Update/ack
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(53) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_t_read_data0_179_delayed_1_0_198_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_t_read_data0_179_delayed_1_0_198_inst_ack_1, ack => accessMem_v_CP_553_elements(53)); -- 
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	21 
    -- CP-element group 54: 	33 
    -- CP-element group 54: 	45 
    -- CP-element group 54: 	49 
    -- CP-element group 54: 	53 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	56 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 assign_stmt_152_to_assign_stmt_224/CONCAT_u32_u64_209_sample_start_
      -- CP-element group 54: 	 assign_stmt_152_to_assign_stmt_224/CONCAT_u32_u64_209_Sample/$entry
      -- CP-element group 54: 	 assign_stmt_152_to_assign_stmt_224/CONCAT_u32_u64_209_Sample/rr
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(54) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:CONCAT_u32_u64_209_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(54), ack => CONCAT_u32_u64_209_inst_req_0); -- 
    accessMem_v_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(21) & accessMem_v_CP_553_elements(33) & accessMem_v_CP_553_elements(45) & accessMem_v_CP_553_elements(49) & accessMem_v_CP_553_elements(53) & accessMem_v_CP_553_elements(56);
      gj_accessMem_v_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	57 
    -- CP-element group 55: 	68 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 assign_stmt_152_to_assign_stmt_224/CONCAT_u32_u64_209_update_start_
      -- CP-element group 55: 	 assign_stmt_152_to_assign_stmt_224/CONCAT_u32_u64_209_Update/$entry
      -- CP-element group 55: 	 assign_stmt_152_to_assign_stmt_224/CONCAT_u32_u64_209_Update/cr
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(55) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:CONCAT_u32_u64_209_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(55), ack => CONCAT_u32_u64_209_inst_req_1); -- 
    accessMem_v_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(57) & accessMem_v_CP_553_elements(68);
      gj_accessMem_v_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	19 
    -- CP-element group 56: 	31 
    -- CP-element group 56: 	43 
    -- CP-element group 56: 	47 
    -- CP-element group 56: 	51 
    -- CP-element group 56: 	54 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 assign_stmt_152_to_assign_stmt_224/CONCAT_u32_u64_209_sample_completed_
      -- CP-element group 56: 	 assign_stmt_152_to_assign_stmt_224/CONCAT_u32_u64_209_Sample/$exit
      -- CP-element group 56: 	 assign_stmt_152_to_assign_stmt_224/CONCAT_u32_u64_209_Sample/ra
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(56) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:CONCAT_u32_u64_209_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_209_inst_ack_0, ack => accessMem_v_CP_553_elements(56)); -- 
    -- CP-element group 57:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	66 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	55 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 assign_stmt_152_to_assign_stmt_224/CONCAT_u32_u64_209_update_completed_
      -- CP-element group 57: 	 assign_stmt_152_to_assign_stmt_224/CONCAT_u32_u64_209_Update/$exit
      -- CP-element group 57: 	 assign_stmt_152_to_assign_stmt_224/CONCAT_u32_u64_209_Update/ca
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(57) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:CONCAT_u32_u64_209_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_209_inst_ack_1, ack => accessMem_v_CP_553_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	1 
    -- CP-element group 58: 	70 
    -- CP-element group 58: 	71 
    -- CP-element group 58: 	72 
    -- CP-element group 58: 	73 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_sample_start_
      -- CP-element group 58: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_Sample/$entry
      -- CP-element group 58: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_Sample/array_obj_ref_213_Split/$entry
      -- CP-element group 58: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_Sample/array_obj_ref_213_Split/$exit
      -- CP-element group 58: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_Sample/array_obj_ref_213_Split/split_req
      -- CP-element group 58: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_Sample/array_obj_ref_213_Split/split_ack
      -- CP-element group 58: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_Sample/word_access_start/$entry
      -- CP-element group 58: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_Sample/word_access_start/word_0/$entry
      -- CP-element group 58: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(58) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:array_obj_ref_213_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(58), ack => array_obj_ref_213_store_0_req_0); -- 
    accessMem_v_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 14,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(1) & accessMem_v_CP_553_elements(70) & accessMem_v_CP_553_elements(71) & accessMem_v_CP_553_elements(72) & accessMem_v_CP_553_elements(73) & accessMem_v_CP_553_elements(60);
      gj_accessMem_v_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (5) 
      -- CP-element group 59: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_update_start_
      -- CP-element group 59: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_Update/$entry
      -- CP-element group 59: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_Update/word_access_complete/$entry
      -- CP-element group 59: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_Update/word_access_complete/word_0/$entry
      -- CP-element group 59: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(59) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:array_obj_ref_213_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(59), ack => array_obj_ref_213_store_0_req_1); -- 
    accessMem_v_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMem_v_CP_553_elements(61);
      gj_accessMem_v_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	74 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	2 
    -- CP-element group 60: 	3 
    -- CP-element group 60: 	4 
    -- CP-element group 60: 	6 
    -- CP-element group 60: 	18 
    -- CP-element group 60: 	30 
    -- CP-element group 60: 	42 
    -- CP-element group 60: 	58 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_sample_completed_
      -- CP-element group 60: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_Sample/$exit
      -- CP-element group 60: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_Sample/word_access_start/$exit
      -- CP-element group 60: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_Sample/word_access_start/word_0/$exit
      -- CP-element group 60: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_Sample/word_access_start/word_0/ra
      -- CP-element group 60: 	 assign_stmt_152_to_assign_stmt_224/ring_reenable_memory_space_5
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(60) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:array_obj_ref_213_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_213_store_0_ack_0, ack => accessMem_v_CP_553_elements(60)); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	74 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (5) 
      -- CP-element group 61: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_update_completed_
      -- CP-element group 61: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_Update/$exit
      -- CP-element group 61: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_Update/word_access_complete/$exit
      -- CP-element group 61: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_Update/word_access_complete/word_0/$exit
      -- CP-element group 61: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_213_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(61) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:array_obj_ref_213_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_213_store_0_ack_1, ack => accessMem_v_CP_553_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	1 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_218_sample_start_
      -- CP-element group 62: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_218_Sample/$entry
      -- CP-element group 62: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_218_Sample/req
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(62) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_read_write_bar_189_delayed_7_0_216_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(62), ack => W_read_write_bar_189_delayed_7_0_216_inst_req_0); -- 
    accessMem_v_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 14,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(1) & accessMem_v_CP_553_elements(64);
      gj_accessMem_v_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: 	68 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_218_update_start_
      -- CP-element group 63: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_218_Update/$entry
      -- CP-element group 63: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_218_Update/req
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(63) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_read_write_bar_189_delayed_7_0_216_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(63), ack => W_read_write_bar_189_delayed_7_0_216_inst_req_1); -- 
    accessMem_v_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(65) & accessMem_v_CP_553_elements(68);
      gj_accessMem_v_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	2 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_218_sample_completed_
      -- CP-element group 64: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_218_Sample/$exit
      -- CP-element group 64: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_218_Sample/ack
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(64) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_read_write_bar_189_delayed_7_0_216_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_189_delayed_7_0_216_inst_ack_0, ack => accessMem_v_CP_553_elements(64)); -- 
    -- CP-element group 65:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65: marked-successors 
    -- CP-element group 65: 	63 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_218_update_completed_
      -- CP-element group 65: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_218_Update/$exit
      -- CP-element group 65: 	 assign_stmt_152_to_assign_stmt_224/assign_stmt_218_Update/ack
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(65) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:W_read_write_bar_189_delayed_7_0_216_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_189_delayed_7_0_216_inst_ack_1, ack => accessMem_v_CP_553_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	57 
    -- CP-element group 66: 	65 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	68 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 assign_stmt_152_to_assign_stmt_224/MUX_223_sample_start_
      -- CP-element group 66: 	 assign_stmt_152_to_assign_stmt_224/MUX_223_start/$entry
      -- CP-element group 66: 	 assign_stmt_152_to_assign_stmt_224/MUX_223_start/req
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(66) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:MUX_223_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(66), ack => MUX_223_inst_req_0); -- 
    accessMem_v_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(57) & accessMem_v_CP_553_elements(65) & accessMem_v_CP_553_elements(68);
      gj_accessMem_v_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	5 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 assign_stmt_152_to_assign_stmt_224/MUX_223_update_start_
      -- CP-element group 67: 	 assign_stmt_152_to_assign_stmt_224/MUX_223_complete/$entry
      -- CP-element group 67: 	 assign_stmt_152_to_assign_stmt_224/MUX_223_complete/req
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(67) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:MUX_223_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_v_CP_553_elements(67), ack => MUX_223_inst_req_1); -- 
    accessMem_v_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 14,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(5) & accessMem_v_CP_553_elements(69);
      gj_accessMem_v_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	55 
    -- CP-element group 68: 	63 
    -- CP-element group 68: 	66 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 assign_stmt_152_to_assign_stmt_224/MUX_223_sample_completed_
      -- CP-element group 68: 	 assign_stmt_152_to_assign_stmt_224/MUX_223_start/$exit
      -- CP-element group 68: 	 assign_stmt_152_to_assign_stmt_224/MUX_223_start/ack
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(68) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:MUX_223_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_223_inst_ack_0, ack => accessMem_v_CP_553_elements(68)); -- 
    -- CP-element group 69:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	74 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	67 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 assign_stmt_152_to_assign_stmt_224/MUX_223_update_completed_
      -- CP-element group 69: 	 assign_stmt_152_to_assign_stmt_224/MUX_223_complete/$exit
      -- CP-element group 69: 	 assign_stmt_152_to_assign_stmt_224/MUX_223_complete/ack
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(69) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:MUX_223_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_223_inst_ack_1, ack => accessMem_v_CP_553_elements(69)); -- 
    -- CP-element group 70:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	8 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	58 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_151_array_obj_ref_213_delay
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(70)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(70)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(70) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accessMem_v_CP_553_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => accessMem_v_CP_553_elements(8), ack => accessMem_v_CP_553_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	20 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	58 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_165_array_obj_ref_213_delay
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(71)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(71)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(71) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accessMem_v_CP_553_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => accessMem_v_CP_553_elements(20), ack => accessMem_v_CP_553_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	32 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	58 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_179_array_obj_ref_213_delay
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(72)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(72)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(72) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accessMem_v_CP_553_elements(72) is a control-delay.
    cp_element_72_delay: control_delay_element  generic map(name => " 72_delay", delay_value => 1)  port map(req => accessMem_v_CP_553_elements(32), ack => accessMem_v_CP_553_elements(72), clk => clk, reset =>reset);
    -- CP-element group 73:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	44 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	58 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 assign_stmt_152_to_assign_stmt_224/array_obj_ref_193_array_obj_ref_213_delay
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(73)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(73)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(73) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accessMem_v_CP_553_elements(73) is a control-delay.
    cp_element_73_delay: control_delay_element  generic map(name => " 73_delay", delay_value => 1)  port map(req => accessMem_v_CP_553_elements(44), ack => accessMem_v_CP_553_elements(73), clk => clk, reset =>reset);
    -- CP-element group 74:  join  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	60 
    -- CP-element group 74: 	61 
    -- CP-element group 74: 	69 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	79 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 assign_stmt_152_to_assign_stmt_224/$exit
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(74)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(74)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(74) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_v_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 14,1 => 14,2 => 14);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "accessMem_v_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMem_v_CP_553_elements(60) & accessMem_v_CP_553_elements(61) & accessMem_v_CP_553_elements(69);
      gj_accessMem_v_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_v_CP_553_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  place  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	2 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 read_write_bar_update_enable
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(75)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(75)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(75) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_v_CP_553_elements(75) <= accessMem_v_CP_553_elements(2);
    -- CP-element group 76:  place  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	3 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 addr_update_enable
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(76)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(76)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(76) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_v_CP_553_elements(76) <= accessMem_v_CP_553_elements(3);
    -- CP-element group 77:  place  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	4 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 write_data_update_enable
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(77)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(77)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(77) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_v_CP_553_elements(77) <= accessMem_v_CP_553_elements(4);
    -- CP-element group 78:  place  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	5 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 read_datal_update_enable
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(78)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(78)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(78) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 79:  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	74 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 $exit
      -- 
    -- logger for CP element group accessMem_v_CP_553_elements(79)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_v_CP_553_elements(79)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem_v:CP:accessMem_v_CP_553_elements(79) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_v_CP_553_elements(79) <= accessMem_v_CP_553_elements(74);
    --  hookup: inputs to control-path 
    accessMem_v_CP_553_elements(78) <= read_datal_update_enable;
    -- hookup: output from control-path 
    read_write_bar_update_enable <= accessMem_v_CP_553_elements(75);
    addr_update_enable <= accessMem_v_CP_553_elements(76);
    write_data_update_enable <= accessMem_v_CP_553_elements(77);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u16_u32_205_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_208_wire : std_logic_vector(31 downto 0);
    signal R_addr1_164_resized : std_logic_vector(10 downto 0);
    signal R_addr1_164_scaled : std_logic_vector(10 downto 0);
    signal R_addr2_178_resized : std_logic_vector(10 downto 0);
    signal R_addr2_178_scaled : std_logic_vector(10 downto 0);
    signal R_addr3_192_resized : std_logic_vector(10 downto 0);
    signal R_addr3_192_scaled : std_logic_vector(10 downto 0);
    signal R_addr_150_resized : std_logic_vector(10 downto 0);
    signal R_addr_150_scaled : std_logic_vector(10 downto 0);
    signal R_addr_212_resized : std_logic_vector(10 downto 0);
    signal R_addr_212_scaled : std_logic_vector(10 downto 0);
    signal addr1_158 : std_logic_vector(11 downto 0);
    signal addr2_172 : std_logic_vector(11 downto 0);
    signal addr3_186 : std_logic_vector(11 downto 0);
    signal array_obj_ref_151_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_151_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_151_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_151_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_151_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_151_word_address_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_151_word_offset_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_165_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_165_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_165_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_165_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_165_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_165_word_address_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_165_word_offset_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_179_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_179_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_179_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_179_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_179_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_179_word_address_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_179_word_offset_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_193_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_193_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_193_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_193_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_193_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_193_word_address_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_193_word_offset_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_213_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_213_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_213_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_213_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_213_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_213_word_address_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_213_word_offset_0 : std_logic_vector(10 downto 0);
    signal konst_156_wire_constant : std_logic_vector(11 downto 0);
    signal konst_170_wire_constant : std_logic_vector(11 downto 0);
    signal konst_184_wire_constant : std_logic_vector(11 downto 0);
    signal konst_222_wire_constant : std_logic_vector(63 downto 0);
    signal read_write_bar_146_delayed_1_0_161 : std_logic_vector(0 downto 0);
    signal read_write_bar_157_delayed_1_0_175 : std_logic_vector(0 downto 0);
    signal read_write_bar_168_delayed_1_0_189 : std_logic_vector(0 downto 0);
    signal read_write_bar_173_delayed_6_0_197 : std_logic_vector(0 downto 0);
    signal read_write_bar_189_delayed_7_0_218 : std_logic_vector(0 downto 0);
    signal t_read_data0_152 : std_logic_vector(15 downto 0);
    signal t_read_data0_179_delayed_1_0_200 : std_logic_vector(15 downto 0);
    signal t_read_data1_166 : std_logic_vector(15 downto 0);
    signal t_read_data2_180 : std_logic_vector(15 downto 0);
    signal t_read_data3_194 : std_logic_vector(15 downto 0);
    signal t_read_datal_210 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_151_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_151_resized_base_address <= "00000000000";
    array_obj_ref_151_word_offset_0 <= "00000000000";
    array_obj_ref_165_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_165_resized_base_address <= "00000000000";
    array_obj_ref_165_word_offset_0 <= "00000000000";
    array_obj_ref_179_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_179_resized_base_address <= "00000000000";
    array_obj_ref_179_word_offset_0 <= "00000000000";
    array_obj_ref_193_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_193_resized_base_address <= "00000000000";
    array_obj_ref_193_word_offset_0 <= "00000000000";
    array_obj_ref_213_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_213_resized_base_address <= "00000000000";
    array_obj_ref_213_word_offset_0 <= "00000000000";
    konst_156_wire_constant <= "000000100000";
    konst_170_wire_constant <= "000001000000";
    konst_184_wire_constant <= "000001100000";
    konst_222_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- logger for split-operator MUX_223_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if MUX_223_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:MUX_223_inst:started:   inputs: " & " read_write_bar_189_delayed_7_0_218 = "& Convert_SLV_To_Hex_String(read_write_bar_189_delayed_7_0_218) & " t_read_datal_210 = "& Convert_SLV_To_Hex_String(t_read_datal_210) & " konst_222_wire_constant = "& Convert_SLV_To_Hex_String(konst_222_wire_constant));
          --
        end if; 
        if MUX_223_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:MUX_223_inst:finished:  outputs: " & " read_datal_buffer= "  & Convert_SLV_To_Hex_String(read_datal_buffer));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    MUX_223_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_223_inst_req_0;
      MUX_223_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_223_inst_req_1;
      MUX_223_inst_ack_1<= update_ack(0);
      MUX_223_inst: SelectSplitProtocol generic map(name => "MUX_223_inst", data_width => 64, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => t_read_datal_210, y => konst_222_wire_constant, sel => read_write_bar_189_delayed_7_0_218, z => read_datal_buffer, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator W_read_write_bar_146_delayed_1_0_159_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_read_write_bar_146_delayed_1_0_159_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:W_read_write_bar_146_delayed_1_0_159_inst:started:   inputs: " & " read_write_bar_buffer = "& Convert_SLV_To_Hex_String(read_write_bar_buffer));
          --
        end if; 
        if W_read_write_bar_146_delayed_1_0_159_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:W_read_write_bar_146_delayed_1_0_159_inst:finished:  outputs: " & " read_write_bar_146_delayed_1_0_161= "  & Convert_SLV_To_Hex_String(read_write_bar_146_delayed_1_0_161));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_read_write_bar_146_delayed_1_0_159_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_write_bar_146_delayed_1_0_159_inst_req_0;
      W_read_write_bar_146_delayed_1_0_159_inst_ack_0<= wack(0);
      rreq(0) <= W_read_write_bar_146_delayed_1_0_159_inst_req_1;
      W_read_write_bar_146_delayed_1_0_159_inst_ack_1<= rack(0);
      W_read_write_bar_146_delayed_1_0_159_inst : InterlockBuffer generic map ( -- 
        name => "W_read_write_bar_146_delayed_1_0_159_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_write_bar_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_write_bar_146_delayed_1_0_161,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_read_write_bar_157_delayed_1_0_173_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_read_write_bar_157_delayed_1_0_173_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:W_read_write_bar_157_delayed_1_0_173_inst:started:   inputs: " & " read_write_bar_buffer = "& Convert_SLV_To_Hex_String(read_write_bar_buffer));
          --
        end if; 
        if W_read_write_bar_157_delayed_1_0_173_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:W_read_write_bar_157_delayed_1_0_173_inst:finished:  outputs: " & " read_write_bar_157_delayed_1_0_175= "  & Convert_SLV_To_Hex_String(read_write_bar_157_delayed_1_0_175));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_read_write_bar_157_delayed_1_0_173_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_write_bar_157_delayed_1_0_173_inst_req_0;
      W_read_write_bar_157_delayed_1_0_173_inst_ack_0<= wack(0);
      rreq(0) <= W_read_write_bar_157_delayed_1_0_173_inst_req_1;
      W_read_write_bar_157_delayed_1_0_173_inst_ack_1<= rack(0);
      W_read_write_bar_157_delayed_1_0_173_inst : InterlockBuffer generic map ( -- 
        name => "W_read_write_bar_157_delayed_1_0_173_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_write_bar_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_write_bar_157_delayed_1_0_175,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_read_write_bar_168_delayed_1_0_187_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_read_write_bar_168_delayed_1_0_187_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:W_read_write_bar_168_delayed_1_0_187_inst:started:   inputs: " & " read_write_bar_buffer = "& Convert_SLV_To_Hex_String(read_write_bar_buffer));
          --
        end if; 
        if W_read_write_bar_168_delayed_1_0_187_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:W_read_write_bar_168_delayed_1_0_187_inst:finished:  outputs: " & " read_write_bar_168_delayed_1_0_189= "  & Convert_SLV_To_Hex_String(read_write_bar_168_delayed_1_0_189));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_read_write_bar_168_delayed_1_0_187_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_write_bar_168_delayed_1_0_187_inst_req_0;
      W_read_write_bar_168_delayed_1_0_187_inst_ack_0<= wack(0);
      rreq(0) <= W_read_write_bar_168_delayed_1_0_187_inst_req_1;
      W_read_write_bar_168_delayed_1_0_187_inst_ack_1<= rack(0);
      W_read_write_bar_168_delayed_1_0_187_inst : InterlockBuffer generic map ( -- 
        name => "W_read_write_bar_168_delayed_1_0_187_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_write_bar_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_write_bar_168_delayed_1_0_189,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_read_write_bar_173_delayed_6_0_195_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_read_write_bar_173_delayed_6_0_195_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:W_read_write_bar_173_delayed_6_0_195_inst:started:   inputs: " & " read_write_bar_buffer = "& Convert_SLV_To_Hex_String(read_write_bar_buffer));
          --
        end if; 
        if W_read_write_bar_173_delayed_6_0_195_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:W_read_write_bar_173_delayed_6_0_195_inst:finished:  outputs: " & " read_write_bar_173_delayed_6_0_197= "  & Convert_SLV_To_Hex_String(read_write_bar_173_delayed_6_0_197));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_read_write_bar_173_delayed_6_0_195_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_write_bar_173_delayed_6_0_195_inst_req_0;
      W_read_write_bar_173_delayed_6_0_195_inst_ack_0<= wack(0);
      rreq(0) <= W_read_write_bar_173_delayed_6_0_195_inst_req_1;
      W_read_write_bar_173_delayed_6_0_195_inst_ack_1<= rack(0);
      W_read_write_bar_173_delayed_6_0_195_inst : InterlockBuffer generic map ( -- 
        name => "W_read_write_bar_173_delayed_6_0_195_inst",
        buffer_size => 6,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_write_bar_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_write_bar_173_delayed_6_0_197,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_read_write_bar_189_delayed_7_0_216_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_read_write_bar_189_delayed_7_0_216_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:W_read_write_bar_189_delayed_7_0_216_inst:started:   inputs: " & " read_write_bar_buffer = "& Convert_SLV_To_Hex_String(read_write_bar_buffer));
          --
        end if; 
        if W_read_write_bar_189_delayed_7_0_216_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:W_read_write_bar_189_delayed_7_0_216_inst:finished:  outputs: " & " read_write_bar_189_delayed_7_0_218= "  & Convert_SLV_To_Hex_String(read_write_bar_189_delayed_7_0_218));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_read_write_bar_189_delayed_7_0_216_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_write_bar_189_delayed_7_0_216_inst_req_0;
      W_read_write_bar_189_delayed_7_0_216_inst_ack_0<= wack(0);
      rreq(0) <= W_read_write_bar_189_delayed_7_0_216_inst_req_1;
      W_read_write_bar_189_delayed_7_0_216_inst_ack_1<= rack(0);
      W_read_write_bar_189_delayed_7_0_216_inst : InterlockBuffer generic map ( -- 
        name => "W_read_write_bar_189_delayed_7_0_216_inst",
        buffer_size => 7,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_write_bar_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_write_bar_189_delayed_7_0_218,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_t_read_data0_179_delayed_1_0_198_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_t_read_data0_179_delayed_1_0_198_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:W_t_read_data0_179_delayed_1_0_198_inst:started:   inputs: " & " t_read_data0_152 = "& Convert_SLV_To_Hex_String(t_read_data0_152));
          --
        end if; 
        if W_t_read_data0_179_delayed_1_0_198_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:W_t_read_data0_179_delayed_1_0_198_inst:finished:  outputs: " & " t_read_data0_179_delayed_1_0_200= "  & Convert_SLV_To_Hex_String(t_read_data0_179_delayed_1_0_200));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_t_read_data0_179_delayed_1_0_198_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_t_read_data0_179_delayed_1_0_198_inst_req_0;
      W_t_read_data0_179_delayed_1_0_198_inst_ack_0<= wack(0);
      rreq(0) <= W_t_read_data0_179_delayed_1_0_198_inst_req_1;
      W_t_read_data0_179_delayed_1_0_198_inst_ack_1<= rack(0);
      W_t_read_data0_179_delayed_1_0_198_inst : InterlockBuffer generic map ( -- 
        name => "W_t_read_data0_179_delayed_1_0_198_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => t_read_data0_152,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => t_read_data0_179_delayed_1_0_200,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for operator array_obj_ref_151_addr_0 flow-through 
    process(array_obj_ref_151_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_151_addr_0:flowthrough  inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " array_obj_ref_151_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_151_root_address) & "outputs: " & " array_obj_ref_151_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_151_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_151_addr_0
    process(array_obj_ref_151_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_151_root_address;
      ov(10 downto 0) := iv;
      array_obj_ref_151_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_151_gather_scatter flow-through 
    process(t_read_data0_152) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_151_gather_scatter:flowthrough  inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " array_obj_ref_151_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_151_data_0) & "outputs: " & " t_read_data0_152= "  & Convert_SLV_To_Hex_String(t_read_data0_152));
      --
    end process; 
    -- equivalence array_obj_ref_151_gather_scatter
    process(array_obj_ref_151_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_151_data_0;
      ov(15 downto 0) := iv;
      t_read_data0_152 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_151_index_0_rename flow-through 
    process(R_addr_150_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_151_index_0_rename:flowthrough  inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " R_addr_150_resized = "& Convert_SLV_To_Hex_String(R_addr_150_resized) & "outputs: " & " R_addr_150_scaled= "  & Convert_SLV_To_Hex_String(R_addr_150_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_151_index_0_rename
    process(R_addr_150_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_150_resized;
      ov(10 downto 0) := iv;
      R_addr_150_scaled <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_151_index_0_resize flow-through 
    process(R_addr_150_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_151_index_0_resize:flowthrough  inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " addr_buffer = "& Convert_SLV_To_Hex_String(addr_buffer) & "outputs: " & " R_addr_150_resized= "  & Convert_SLV_To_Hex_String(R_addr_150_resized));
      --
    end process; 
    -- equivalence array_obj_ref_151_index_0_resize
    process(addr_buffer) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_buffer;
      ov := iv(10 downto 0);
      R_addr_150_resized <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_151_index_offset flow-through 
    process(array_obj_ref_151_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_151_index_offset:flowthrough  inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " R_addr_150_scaled = "& Convert_SLV_To_Hex_String(R_addr_150_scaled) & "outputs: " & " array_obj_ref_151_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_151_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_151_index_offset
    process(R_addr_150_scaled) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_150_scaled;
      ov(10 downto 0) := iv;
      array_obj_ref_151_final_offset <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_151_root_address_inst flow-through 
    process(array_obj_ref_151_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_151_root_address_inst:flowthrough  inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " array_obj_ref_151_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_151_final_offset) & "outputs: " & " array_obj_ref_151_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_151_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_151_root_address_inst
    process(array_obj_ref_151_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_151_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_151_root_address <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_165_addr_0 flow-through 
    process(array_obj_ref_165_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_165_addr_0:flowthrough  inputs: " & " read_write_bar_146_delayed_1_0_161 (guard)= " & Convert_SLV_To_String(read_write_bar_146_delayed_1_0_161) & " array_obj_ref_165_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_165_root_address) & "outputs: " & " array_obj_ref_165_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_165_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_165_addr_0
    process(array_obj_ref_165_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_165_root_address;
      ov(10 downto 0) := iv;
      array_obj_ref_165_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_165_gather_scatter flow-through 
    process(t_read_data1_166) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_165_gather_scatter:flowthrough  inputs: " & " read_write_bar_146_delayed_1_0_161 (guard)= " & Convert_SLV_To_String(read_write_bar_146_delayed_1_0_161) & " array_obj_ref_165_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_165_data_0) & "outputs: " & " t_read_data1_166= "  & Convert_SLV_To_Hex_String(t_read_data1_166));
      --
    end process; 
    -- equivalence array_obj_ref_165_gather_scatter
    process(array_obj_ref_165_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_165_data_0;
      ov(15 downto 0) := iv;
      t_read_data1_166 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_165_index_0_rename flow-through 
    process(R_addr1_164_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_165_index_0_rename:flowthrough  inputs: " & " read_write_bar_146_delayed_1_0_161 (guard)= " & Convert_SLV_To_String(read_write_bar_146_delayed_1_0_161) & " R_addr1_164_resized = "& Convert_SLV_To_Hex_String(R_addr1_164_resized) & "outputs: " & " R_addr1_164_scaled= "  & Convert_SLV_To_Hex_String(R_addr1_164_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_165_index_0_rename
    process(R_addr1_164_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr1_164_resized;
      ov(10 downto 0) := iv;
      R_addr1_164_scaled <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_165_index_0_resize flow-through 
    process(R_addr1_164_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_165_index_0_resize:flowthrough  inputs: " & " read_write_bar_146_delayed_1_0_161 (guard)= " & Convert_SLV_To_String(read_write_bar_146_delayed_1_0_161) & " addr1_158 = "& Convert_SLV_To_Hex_String(addr1_158) & "outputs: " & " R_addr1_164_resized= "  & Convert_SLV_To_Hex_String(R_addr1_164_resized));
      --
    end process; 
    -- equivalence array_obj_ref_165_index_0_resize
    process(addr1_158) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr1_158;
      ov := iv(10 downto 0);
      R_addr1_164_resized <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_165_index_offset flow-through 
    process(array_obj_ref_165_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_165_index_offset:flowthrough  inputs: " & " read_write_bar_146_delayed_1_0_161 (guard)= " & Convert_SLV_To_String(read_write_bar_146_delayed_1_0_161) & " R_addr1_164_scaled = "& Convert_SLV_To_Hex_String(R_addr1_164_scaled) & "outputs: " & " array_obj_ref_165_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_165_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_165_index_offset
    process(R_addr1_164_scaled) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr1_164_scaled;
      ov(10 downto 0) := iv;
      array_obj_ref_165_final_offset <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_165_root_address_inst flow-through 
    process(array_obj_ref_165_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_165_root_address_inst:flowthrough  inputs: " & " read_write_bar_146_delayed_1_0_161 (guard)= " & Convert_SLV_To_String(read_write_bar_146_delayed_1_0_161) & " array_obj_ref_165_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_165_final_offset) & "outputs: " & " array_obj_ref_165_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_165_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_165_root_address_inst
    process(array_obj_ref_165_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_165_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_165_root_address <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_179_addr_0 flow-through 
    process(array_obj_ref_179_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_179_addr_0:flowthrough  inputs: " & " read_write_bar_157_delayed_1_0_175 (guard)= " & Convert_SLV_To_String(read_write_bar_157_delayed_1_0_175) & " array_obj_ref_179_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_179_root_address) & "outputs: " & " array_obj_ref_179_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_179_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_179_addr_0
    process(array_obj_ref_179_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_179_root_address;
      ov(10 downto 0) := iv;
      array_obj_ref_179_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_179_gather_scatter flow-through 
    process(t_read_data2_180) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_179_gather_scatter:flowthrough  inputs: " & " read_write_bar_157_delayed_1_0_175 (guard)= " & Convert_SLV_To_String(read_write_bar_157_delayed_1_0_175) & " array_obj_ref_179_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_179_data_0) & "outputs: " & " t_read_data2_180= "  & Convert_SLV_To_Hex_String(t_read_data2_180));
      --
    end process; 
    -- equivalence array_obj_ref_179_gather_scatter
    process(array_obj_ref_179_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_179_data_0;
      ov(15 downto 0) := iv;
      t_read_data2_180 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_179_index_0_rename flow-through 
    process(R_addr2_178_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_179_index_0_rename:flowthrough  inputs: " & " read_write_bar_157_delayed_1_0_175 (guard)= " & Convert_SLV_To_String(read_write_bar_157_delayed_1_0_175) & " R_addr2_178_resized = "& Convert_SLV_To_Hex_String(R_addr2_178_resized) & "outputs: " & " R_addr2_178_scaled= "  & Convert_SLV_To_Hex_String(R_addr2_178_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_179_index_0_rename
    process(R_addr2_178_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr2_178_resized;
      ov(10 downto 0) := iv;
      R_addr2_178_scaled <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_179_index_0_resize flow-through 
    process(R_addr2_178_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_179_index_0_resize:flowthrough  inputs: " & " read_write_bar_157_delayed_1_0_175 (guard)= " & Convert_SLV_To_String(read_write_bar_157_delayed_1_0_175) & " addr2_172 = "& Convert_SLV_To_Hex_String(addr2_172) & "outputs: " & " R_addr2_178_resized= "  & Convert_SLV_To_Hex_String(R_addr2_178_resized));
      --
    end process; 
    -- equivalence array_obj_ref_179_index_0_resize
    process(addr2_172) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr2_172;
      ov := iv(10 downto 0);
      R_addr2_178_resized <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_179_index_offset flow-through 
    process(array_obj_ref_179_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_179_index_offset:flowthrough  inputs: " & " read_write_bar_157_delayed_1_0_175 (guard)= " & Convert_SLV_To_String(read_write_bar_157_delayed_1_0_175) & " R_addr2_178_scaled = "& Convert_SLV_To_Hex_String(R_addr2_178_scaled) & "outputs: " & " array_obj_ref_179_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_179_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_179_index_offset
    process(R_addr2_178_scaled) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr2_178_scaled;
      ov(10 downto 0) := iv;
      array_obj_ref_179_final_offset <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_179_root_address_inst flow-through 
    process(array_obj_ref_179_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_179_root_address_inst:flowthrough  inputs: " & " read_write_bar_157_delayed_1_0_175 (guard)= " & Convert_SLV_To_String(read_write_bar_157_delayed_1_0_175) & " array_obj_ref_179_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_179_final_offset) & "outputs: " & " array_obj_ref_179_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_179_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_179_root_address_inst
    process(array_obj_ref_179_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_179_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_179_root_address <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_193_addr_0 flow-through 
    process(array_obj_ref_193_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_193_addr_0:flowthrough  inputs: " & " read_write_bar_168_delayed_1_0_189 (guard)= " & Convert_SLV_To_String(read_write_bar_168_delayed_1_0_189) & " array_obj_ref_193_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_193_root_address) & "outputs: " & " array_obj_ref_193_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_193_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_193_addr_0
    process(array_obj_ref_193_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_193_root_address;
      ov(10 downto 0) := iv;
      array_obj_ref_193_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_193_gather_scatter flow-through 
    process(t_read_data3_194) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_193_gather_scatter:flowthrough  inputs: " & " read_write_bar_168_delayed_1_0_189 (guard)= " & Convert_SLV_To_String(read_write_bar_168_delayed_1_0_189) & " array_obj_ref_193_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_193_data_0) & "outputs: " & " t_read_data3_194= "  & Convert_SLV_To_Hex_String(t_read_data3_194));
      --
    end process; 
    -- equivalence array_obj_ref_193_gather_scatter
    process(array_obj_ref_193_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_193_data_0;
      ov(15 downto 0) := iv;
      t_read_data3_194 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_193_index_0_rename flow-through 
    process(R_addr3_192_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_193_index_0_rename:flowthrough  inputs: " & " read_write_bar_168_delayed_1_0_189 (guard)= " & Convert_SLV_To_String(read_write_bar_168_delayed_1_0_189) & " R_addr3_192_resized = "& Convert_SLV_To_Hex_String(R_addr3_192_resized) & "outputs: " & " R_addr3_192_scaled= "  & Convert_SLV_To_Hex_String(R_addr3_192_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_193_index_0_rename
    process(R_addr3_192_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr3_192_resized;
      ov(10 downto 0) := iv;
      R_addr3_192_scaled <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_193_index_0_resize flow-through 
    process(R_addr3_192_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_193_index_0_resize:flowthrough  inputs: " & " read_write_bar_168_delayed_1_0_189 (guard)= " & Convert_SLV_To_String(read_write_bar_168_delayed_1_0_189) & " addr3_186 = "& Convert_SLV_To_Hex_String(addr3_186) & "outputs: " & " R_addr3_192_resized= "  & Convert_SLV_To_Hex_String(R_addr3_192_resized));
      --
    end process; 
    -- equivalence array_obj_ref_193_index_0_resize
    process(addr3_186) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr3_186;
      ov := iv(10 downto 0);
      R_addr3_192_resized <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_193_index_offset flow-through 
    process(array_obj_ref_193_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_193_index_offset:flowthrough  inputs: " & " read_write_bar_168_delayed_1_0_189 (guard)= " & Convert_SLV_To_String(read_write_bar_168_delayed_1_0_189) & " R_addr3_192_scaled = "& Convert_SLV_To_Hex_String(R_addr3_192_scaled) & "outputs: " & " array_obj_ref_193_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_193_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_193_index_offset
    process(R_addr3_192_scaled) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr3_192_scaled;
      ov(10 downto 0) := iv;
      array_obj_ref_193_final_offset <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_193_root_address_inst flow-through 
    process(array_obj_ref_193_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_193_root_address_inst:flowthrough  inputs: " & " read_write_bar_168_delayed_1_0_189 (guard)= " & Convert_SLV_To_String(read_write_bar_168_delayed_1_0_189) & " array_obj_ref_193_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_193_final_offset) & "outputs: " & " array_obj_ref_193_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_193_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_193_root_address_inst
    process(array_obj_ref_193_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_193_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_193_root_address <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_213_addr_0 flow-through 
    process(array_obj_ref_213_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_213_addr_0:flowthrough  inputs: " & " read_write_bar_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_buffer) & " array_obj_ref_213_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_213_root_address) & "outputs: " & " array_obj_ref_213_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_213_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_213_addr_0
    process(array_obj_ref_213_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_213_root_address;
      ov(10 downto 0) := iv;
      array_obj_ref_213_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_213_gather_scatter flow-through 
    process(array_obj_ref_213_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_213_gather_scatter:flowthrough  inputs: " & " read_write_bar_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_buffer) & " write_data_buffer = "& Convert_SLV_To_Hex_String(write_data_buffer) & "outputs: " & " array_obj_ref_213_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_213_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_213_gather_scatter
    process(write_data_buffer) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := write_data_buffer;
      ov(15 downto 0) := iv;
      array_obj_ref_213_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_213_index_0_rename flow-through 
    process(R_addr_212_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_213_index_0_rename:flowthrough  inputs: " & " read_write_bar_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_buffer) & " R_addr_212_resized = "& Convert_SLV_To_Hex_String(R_addr_212_resized) & "outputs: " & " R_addr_212_scaled= "  & Convert_SLV_To_Hex_String(R_addr_212_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_213_index_0_rename
    process(R_addr_212_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_212_resized;
      ov(10 downto 0) := iv;
      R_addr_212_scaled <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_213_index_0_resize flow-through 
    process(R_addr_212_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_213_index_0_resize:flowthrough  inputs: " & " read_write_bar_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_buffer) & " addr_buffer = "& Convert_SLV_To_Hex_String(addr_buffer) & "outputs: " & " R_addr_212_resized= "  & Convert_SLV_To_Hex_String(R_addr_212_resized));
      --
    end process; 
    -- equivalence array_obj_ref_213_index_0_resize
    process(addr_buffer) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_buffer;
      ov := iv(10 downto 0);
      R_addr_212_resized <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_213_index_offset flow-through 
    process(array_obj_ref_213_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_213_index_offset:flowthrough  inputs: " & " read_write_bar_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_buffer) & " R_addr_212_scaled = "& Convert_SLV_To_Hex_String(R_addr_212_scaled) & "outputs: " & " array_obj_ref_213_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_213_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_213_index_offset
    process(R_addr_212_scaled) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_212_scaled;
      ov(10 downto 0) := iv;
      array_obj_ref_213_final_offset <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_213_root_address_inst flow-through 
    process(array_obj_ref_213_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_213_root_address_inst:flowthrough  inputs: " & " read_write_bar_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_buffer) & " array_obj_ref_213_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_213_final_offset) & "outputs: " & " array_obj_ref_213_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_213_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_213_root_address_inst
    process(array_obj_ref_213_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_213_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_213_root_address <= ov(10 downto 0);
      --
    end process;
    -- logger for split-operator ADD_u12_u12_157_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_157_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:ADD_u12_u12_157_inst:started:   inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " addr_buffer = "& Convert_SLV_To_Hex_String(addr_buffer) & " konst_156_wire_constant = "& Convert_SLV_To_Hex_String(konst_156_wire_constant));
          --
        end if; 
        if ADD_u12_u12_157_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:ADD_u12_u12_157_inst:finished:  outputs: " & " addr1_158= "  & Convert_SLV_To_Hex_String(addr1_158));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (0) : ADD_u12_u12_157_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= addr_buffer;
      addr1_158 <= data_out(11 downto 0);
      guard_vector(0)  <= read_write_bar_buffer(0);
      reqL_unguarded(0) <= ADD_u12_u12_157_inst_req_0;
      ADD_u12_u12_157_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_157_inst_req_1;
      ADD_u12_u12_157_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000000100000",
          constant_width => 12,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- logger for split-operator ADD_u12_u12_171_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_171_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:ADD_u12_u12_171_inst:started:   inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " addr_buffer = "& Convert_SLV_To_Hex_String(addr_buffer) & " konst_170_wire_constant = "& Convert_SLV_To_Hex_String(konst_170_wire_constant));
          --
        end if; 
        if ADD_u12_u12_171_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:ADD_u12_u12_171_inst:finished:  outputs: " & " addr2_172= "  & Convert_SLV_To_Hex_String(addr2_172));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (1) : ADD_u12_u12_171_inst 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= addr_buffer;
      addr2_172 <= data_out(11 downto 0);
      guard_vector(0)  <= read_write_bar_buffer(0);
      reqL_unguarded(0) <= ADD_u12_u12_171_inst_req_0;
      ADD_u12_u12_171_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_171_inst_req_1;
      ADD_u12_u12_171_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000001000000",
          constant_width => 12,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- logger for split-operator ADD_u12_u12_185_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_185_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:ADD_u12_u12_185_inst:started:   inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " addr_buffer = "& Convert_SLV_To_Hex_String(addr_buffer) & " konst_184_wire_constant = "& Convert_SLV_To_Hex_String(konst_184_wire_constant));
          --
        end if; 
        if ADD_u12_u12_185_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:ADD_u12_u12_185_inst:finished:  outputs: " & " addr3_186= "  & Convert_SLV_To_Hex_String(addr3_186));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (2) : ADD_u12_u12_185_inst 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= addr_buffer;
      addr3_186 <= data_out(11 downto 0);
      guard_vector(0)  <= read_write_bar_buffer(0);
      reqL_unguarded(0) <= ADD_u12_u12_185_inst_req_0;
      ADD_u12_u12_185_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_185_inst_req_1;
      ADD_u12_u12_185_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_2_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000001100000",
          constant_width => 12,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- logger for split-operator CONCAT_u16_u32_205_inst flow-through 
    process(CONCAT_u16_u32_205_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:CONCAT_u16_u32_205_inst:flowthrough inputs: " & " read_write_bar_173_delayed_6_0_197 (guard)= " & Convert_SLV_To_String(read_write_bar_173_delayed_6_0_197) & " t_read_data3_194 = "& Convert_SLV_To_Hex_String(t_read_data3_194) & " t_read_data2_180 = "& Convert_SLV_To_Hex_String(t_read_data2_180) & " outputs:" & " CONCAT_u16_u32_205_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u16_u32_205_wire));
      --
    end process; 
    -- binary operator CONCAT_u16_u32_205_inst
    process(t_read_data3_194, t_read_data2_180) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(t_read_data3_194, t_read_data2_180, tmp_var);
      CONCAT_u16_u32_205_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u16_u32_208_inst flow-through 
    process(CONCAT_u16_u32_208_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:CONCAT_u16_u32_208_inst:flowthrough inputs: " & " read_write_bar_173_delayed_6_0_197 (guard)= " & Convert_SLV_To_String(read_write_bar_173_delayed_6_0_197) & " t_read_data1_166 = "& Convert_SLV_To_Hex_String(t_read_data1_166) & " t_read_data0_179_delayed_1_0_200 = "& Convert_SLV_To_Hex_String(t_read_data0_179_delayed_1_0_200) & " outputs:" & " CONCAT_u16_u32_208_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u16_u32_208_wire));
      --
    end process; 
    -- binary operator CONCAT_u16_u32_208_inst
    process(t_read_data1_166, t_read_data0_179_delayed_1_0_200) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(t_read_data1_166, t_read_data0_179_delayed_1_0_200, tmp_var);
      CONCAT_u16_u32_208_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u32_u64_209_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if CONCAT_u32_u64_209_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:CONCAT_u32_u64_209_inst:started:   inputs: " & " read_write_bar_173_delayed_6_0_197 (guard)= " & Convert_SLV_To_String(read_write_bar_173_delayed_6_0_197) & " CONCAT_u16_u32_205_wire = "& Convert_SLV_To_Hex_String(CONCAT_u16_u32_205_wire) & " CONCAT_u16_u32_208_wire = "& Convert_SLV_To_Hex_String(CONCAT_u16_u32_208_wire));
          --
        end if; 
        if CONCAT_u32_u64_209_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:CONCAT_u32_u64_209_inst:finished:  outputs: " & " t_read_datal_210= "  & Convert_SLV_To_Hex_String(t_read_datal_210));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (5) : CONCAT_u32_u64_209_inst 
    ApConcat_group_5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_205_wire & CONCAT_u16_u32_208_wire;
      t_read_datal_210 <= data_out(63 downto 0);
      guard_vector(0)  <= read_write_bar_173_delayed_6_0_197(0);
      reqL_unguarded(0) <= CONCAT_u32_u64_209_inst_req_0;
      CONCAT_u32_u64_209_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_209_inst_req_1;
      CONCAT_u32_u64_209_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_5_gI: SplitGuardInterface generic map(name => "ApConcat_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- logger for split-operator array_obj_ref_151_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_151_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_151_load_0:started:   inputs: " & " read_write_bar_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_buffer) & " array_obj_ref_151_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_151_word_address_0));
          --
        end if; 
        if array_obj_ref_151_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_151_load_0:finished:  outputs: " & " array_obj_ref_151_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_151_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_165_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_165_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_165_load_0:started:   inputs: " & " read_write_bar_146_delayed_1_0_161 (guard)= " & Convert_SLV_To_String(read_write_bar_146_delayed_1_0_161) & " array_obj_ref_165_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_165_word_address_0));
          --
        end if; 
        if array_obj_ref_165_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_165_load_0:finished:  outputs: " & " array_obj_ref_165_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_165_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_179_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_179_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_179_load_0:started:   inputs: " & " read_write_bar_157_delayed_1_0_175 (guard)= " & Convert_SLV_To_String(read_write_bar_157_delayed_1_0_175) & " array_obj_ref_179_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_179_word_address_0));
          --
        end if; 
        if array_obj_ref_179_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_179_load_0:finished:  outputs: " & " array_obj_ref_179_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_179_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_193_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_193_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_193_load_0:started:   inputs: " & " read_write_bar_168_delayed_1_0_189 (guard)= " & Convert_SLV_To_String(read_write_bar_168_delayed_1_0_189) & " array_obj_ref_193_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_193_word_address_0));
          --
        end if; 
        if array_obj_ref_193_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_193_load_0:finished:  outputs: " & " array_obj_ref_193_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_193_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (0) : array_obj_ref_151_load_0 array_obj_ref_165_load_0 array_obj_ref_179_load_0 array_obj_ref_193_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(43 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => true, 1 => true, 2 => true, 3 => true);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 5, 1 => 5, 2 => 5, 3 => 5);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_151_load_0_req_0,
        array_obj_ref_151_load_0_ack_0,
        array_obj_ref_151_load_0_req_1,
        array_obj_ref_151_load_0_ack_1,
        "array_obj_ref_151_load_0",
        "memory_space_5" ,
        array_obj_ref_151_data_0,
        array_obj_ref_151_word_address_0,
        "array_obj_ref_151_data_0",
        "array_obj_ref_151_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_165_load_0_req_0,
        array_obj_ref_165_load_0_ack_0,
        array_obj_ref_165_load_0_req_1,
        array_obj_ref_165_load_0_ack_1,
        "array_obj_ref_165_load_0",
        "memory_space_5" ,
        array_obj_ref_165_data_0,
        array_obj_ref_165_word_address_0,
        "array_obj_ref_165_data_0",
        "array_obj_ref_165_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_179_load_0_req_0,
        array_obj_ref_179_load_0_ack_0,
        array_obj_ref_179_load_0_req_1,
        array_obj_ref_179_load_0_ack_1,
        "array_obj_ref_179_load_0",
        "memory_space_5" ,
        array_obj_ref_179_data_0,
        array_obj_ref_179_word_address_0,
        "array_obj_ref_179_data_0",
        "array_obj_ref_179_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_193_load_0_req_0,
        array_obj_ref_193_load_0_ack_0,
        array_obj_ref_193_load_0_req_1,
        array_obj_ref_193_load_0_ack_1,
        "array_obj_ref_193_load_0",
        "memory_space_5" ,
        array_obj_ref_193_data_0,
        array_obj_ref_193_word_address_0,
        "array_obj_ref_193_data_0",
        "array_obj_ref_193_word_address_0" -- 
      );
      reqL_unguarded(3) <= array_obj_ref_151_load_0_req_0;
      reqL_unguarded(2) <= array_obj_ref_165_load_0_req_0;
      reqL_unguarded(1) <= array_obj_ref_179_load_0_req_0;
      reqL_unguarded(0) <= array_obj_ref_193_load_0_req_0;
      array_obj_ref_151_load_0_ack_0 <= ackL_unguarded(3);
      array_obj_ref_165_load_0_ack_0 <= ackL_unguarded(2);
      array_obj_ref_179_load_0_ack_0 <= ackL_unguarded(1);
      array_obj_ref_193_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= array_obj_ref_151_load_0_req_1;
      reqR_unguarded(2) <= array_obj_ref_165_load_0_req_1;
      reqR_unguarded(1) <= array_obj_ref_179_load_0_req_1;
      reqR_unguarded(0) <= array_obj_ref_193_load_0_req_1;
      array_obj_ref_151_load_0_ack_1 <= ackR_unguarded(3);
      array_obj_ref_165_load_0_ack_1 <= ackR_unguarded(2);
      array_obj_ref_179_load_0_ack_1 <= ackR_unguarded(1);
      array_obj_ref_193_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_write_bar_168_delayed_1_0_189(0);
      guard_vector(1)  <= read_write_bar_157_delayed_1_0_175(0);
      guard_vector(2)  <= read_write_bar_146_delayed_1_0_161(0);
      guard_vector(3)  <= read_write_bar_buffer(0);
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_151_word_address_0 & array_obj_ref_165_word_address_0 & array_obj_ref_179_word_address_0 & array_obj_ref_193_word_address_0;
      array_obj_ref_151_data_0 <= data_out(63 downto 48);
      array_obj_ref_165_data_0 <= data_out(47 downto 32);
      array_obj_ref_179_data_0 <= data_out(31 downto 16);
      array_obj_ref_193_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 11,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(10 downto 0),
          mtag => memory_space_5_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(15 downto 0),
          mtag => memory_space_5_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logger for split-operator array_obj_ref_213_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_213_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_213_store_0:started:   inputs: " & " read_write_bar_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_buffer) & " array_obj_ref_213_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_213_word_address_0) & " array_obj_ref_213_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_213_data_0));
          --
        end if; 
        if array_obj_ref_213_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem_v:DP:array_obj_ref_213_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_213_store_0_req_0,
      array_obj_ref_213_store_0_ack_0,
      array_obj_ref_213_store_0_req_1,
      array_obj_ref_213_store_0_ack_1,
      "array_obj_ref_213_store_0",
      "memory_space_5" ,
      array_obj_ref_213_data_0,
      array_obj_ref_213_word_address_0,
      "array_obj_ref_213_data_0",
      "array_obj_ref_213_word_address_0" -- 
    );
    -- shared store operator group (0) : array_obj_ref_213_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_213_store_0_req_0;
      array_obj_ref_213_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_213_store_0_req_1;
      array_obj_ref_213_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_write_bar_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_213_word_address_0;
      data_in <= array_obj_ref_213_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 11,
        data_width => 16,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(10 downto 0),
          mdata => memory_space_5_sr_data(15 downto 0),
          mtag => memory_space_5_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end accessMem_v_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity initial is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(11 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(11 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    accessMem_call_reqs : out  std_logic_vector(0 downto 0);
    accessMem_call_acks : in   std_logic_vector(0 downto 0);
    accessMem_call_data : out  std_logic_vector(28 downto 0);
    accessMem_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMem_return_reqs : out  std_logic_vector(0 downto 0);
    accessMem_return_acks : in   std_logic_vector(0 downto 0);
    accessMem_return_data : in   std_logic_vector(63 downto 0);
    accessMem_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity initial;
architecture initial_arch of initial is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal initial_CP_1047_start: Boolean;
  signal initial_CP_1047_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(11 downto 0);
      write_data : in  std_logic_vector(15 downto 0);
      read_datal : out  std_logic_vector(63 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal STORE_ZJ_241_store_0_ack_1 : boolean;
  signal do_while_stmt_247_branch_req_0 : boolean;
  signal STORE_ZJ_241_store_0_req_0 : boolean;
  signal phi_stmt_249_req_1 : boolean;
  signal STORE_ZJ_230_store_0_ack_1 : boolean;
  signal STORE_ZJ_241_store_0_req_1 : boolean;
  signal phi_stmt_249_req_0 : boolean;
  signal NI_280_253_buf_req_0 : boolean;
  signal STORE_ZJ_241_store_0_ack_0 : boolean;
  signal STORE_ZJ_230_store_0_req_0 : boolean;
  signal MUL_u12_u12_244_inst_req_0 : boolean;
  signal MUL_u12_u12_244_inst_ack_0 : boolean;
  signal STORE_ZJ_230_store_0_req_1 : boolean;
  signal NI_280_253_buf_ack_0 : boolean;
  signal NI_280_253_buf_req_1 : boolean;
  signal phi_stmt_249_ack_0 : boolean;
  signal MUL_u12_u12_244_inst_req_1 : boolean;
  signal MUL_u12_u12_244_inst_ack_1 : boolean;
  signal STORE_ZJ_230_store_0_ack_0 : boolean;
  signal W_I_230_delayed_4_0_259_inst_req_0 : boolean;
  signal W_I_230_delayed_4_0_259_inst_ack_0 : boolean;
  signal W_I_230_delayed_4_0_259_inst_req_1 : boolean;
  signal W_I_230_delayed_4_0_259_inst_ack_1 : boolean;
  signal NI_280_253_buf_ack_1 : boolean;
  signal type_cast_257_inst_req_0 : boolean;
  signal type_cast_257_inst_ack_0 : boolean;
  signal type_cast_257_inst_req_1 : boolean;
  signal type_cast_257_inst_ack_1 : boolean;
  signal LOAD_ZJ_263_load_0_req_0 : boolean;
  signal LOAD_ZJ_263_load_0_ack_0 : boolean;
  signal LOAD_ZJ_263_load_0_req_1 : boolean;
  signal LOAD_ZJ_263_load_0_ack_1 : boolean;
  signal type_cast_266_inst_req_0 : boolean;
  signal type_cast_266_inst_ack_0 : boolean;
  signal type_cast_266_inst_req_1 : boolean;
  signal type_cast_266_inst_ack_1 : boolean;
  signal W_wdata_236_delayed_4_0_268_inst_req_0 : boolean;
  signal W_wdata_236_delayed_4_0_268_inst_ack_0 : boolean;
  signal W_wdata_236_delayed_4_0_268_inst_req_1 : boolean;
  signal W_wdata_236_delayed_4_0_268_inst_ack_1 : boolean;
  signal call_stmt_275_call_req_0 : boolean;
  signal call_stmt_275_call_ack_0 : boolean;
  signal call_stmt_275_call_req_1 : boolean;
  signal call_stmt_275_call_ack_1 : boolean;
  signal ADD_u12_u12_279_inst_req_0 : boolean;
  signal ADD_u12_u12_279_inst_ack_0 : boolean;
  signal ADD_u12_u12_279_inst_req_1 : boolean;
  signal ADD_u12_u12_279_inst_ack_1 : boolean;
  signal do_while_stmt_247_branch_ack_0 : boolean;
  signal do_while_stmt_247_branch_ack_1 : boolean;
  signal ADD_u12_u12_289_inst_req_0 : boolean;
  signal ADD_u12_u12_289_inst_ack_0 : boolean;
  signal ADD_u12_u12_289_inst_req_1 : boolean;
  signal ADD_u12_u12_289_inst_ack_1 : boolean;
  signal do_while_stmt_302_branch_ack_1 : boolean;
  signal if_stmt_291_branch_req_0 : boolean;
  signal do_while_stmt_302_branch_ack_0 : boolean;
  signal if_stmt_291_branch_ack_1 : boolean;
  signal if_stmt_291_branch_ack_0 : boolean;
  signal phi_stmt_235_req_0 : boolean;
  signal YI_290_239_buf_req_0 : boolean;
  signal YI_290_239_buf_ack_0 : boolean;
  signal YI_290_239_buf_req_1 : boolean;
  signal YI_290_239_buf_ack_1 : boolean;
  signal phi_stmt_235_req_1 : boolean;
  signal phi_stmt_235_ack_0 : boolean;
  signal STORE_ZJ_298_store_0_req_0 : boolean;
  signal STORE_ZJ_298_store_0_ack_0 : boolean;
  signal STORE_ZJ_298_store_0_req_1 : boolean;
  signal STORE_ZJ_298_store_0_ack_1 : boolean;
  signal do_while_stmt_302_branch_req_0 : boolean;
  signal phi_stmt_304_req_1 : boolean;
  signal phi_stmt_304_req_0 : boolean;
  signal phi_stmt_304_ack_0 : boolean;
  signal NM_335_308_buf_req_0 : boolean;
  signal NM_335_308_buf_ack_0 : boolean;
  signal NM_335_308_buf_req_1 : boolean;
  signal NM_335_308_buf_ack_1 : boolean;
  signal type_cast_312_inst_req_0 : boolean;
  signal type_cast_312_inst_ack_0 : boolean;
  signal type_cast_312_inst_req_1 : boolean;
  signal type_cast_312_inst_ack_1 : boolean;
  signal W_M_279_delayed_4_0_314_inst_req_0 : boolean;
  signal W_M_279_delayed_4_0_314_inst_ack_0 : boolean;
  signal W_M_279_delayed_4_0_314_inst_req_1 : boolean;
  signal W_M_279_delayed_4_0_314_inst_ack_1 : boolean;
  signal LOAD_ZJ_318_load_0_req_0 : boolean;
  signal LOAD_ZJ_318_load_0_ack_0 : boolean;
  signal LOAD_ZJ_318_load_0_req_1 : boolean;
  signal LOAD_ZJ_318_load_0_ack_1 : boolean;
  signal type_cast_321_inst_req_0 : boolean;
  signal type_cast_321_inst_ack_0 : boolean;
  signal type_cast_321_inst_req_1 : boolean;
  signal type_cast_321_inst_ack_1 : boolean;
  signal W_wdata_285_delayed_4_0_323_inst_req_0 : boolean;
  signal W_wdata_285_delayed_4_0_323_inst_ack_0 : boolean;
  signal W_wdata_285_delayed_4_0_323_inst_req_1 : boolean;
  signal W_wdata_285_delayed_4_0_323_inst_ack_1 : boolean;
  signal call_stmt_330_call_req_0 : boolean;
  signal call_stmt_330_call_ack_0 : boolean;
  signal call_stmt_330_call_req_1 : boolean;
  signal call_stmt_330_call_ack_1 : boolean;
  signal ADD_u12_u12_334_inst_req_0 : boolean;
  signal ADD_u12_u12_334_inst_ack_0 : boolean;
  signal ADD_u12_u12_334_inst_req_1 : boolean;
  signal ADD_u12_u12_334_inst_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "initial_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  initial_CP_1047_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "initial_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= initial_CP_1047_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= initial_CP_1047_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= initial_CP_1047_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,initial_CP_1047_start,"initial cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,initial_CP_1047_symbol, "initial cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  initial_CP_1047: Block -- control-path 
    signal initial_CP_1047_elements: BooleanArray(139 downto 0);
    -- 
  begin -- 
    initial_CP_1047_elements(0) <= initial_CP_1047_start;
    initial_CP_1047_symbol <= initial_CP_1047_elements(80);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (18) 
      -- CP-element group 0: 	 assign_stmt_232/STORE_ZJ_230_Sample/STORE_ZJ_230_Split/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_232/STORE_ZJ_230_Update/$entry
      -- CP-element group 0: 	 assign_stmt_232/STORE_ZJ_230_Sample/STORE_ZJ_230_Split/split_ack
      -- CP-element group 0: 	 assign_stmt_232/STORE_ZJ_230_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_232/STORE_ZJ_230_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_232/STORE_ZJ_230_sample_start_
      -- CP-element group 0: 	 assign_stmt_232/STORE_ZJ_230_update_start_
      -- CP-element group 0: 	 assign_stmt_232/$entry
      -- CP-element group 0: 	 assign_stmt_232/STORE_ZJ_230_Sample/STORE_ZJ_230_Split/$exit
      -- CP-element group 0: 	 assign_stmt_232/STORE_ZJ_230_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_232/STORE_ZJ_230_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_232/STORE_ZJ_230_Sample/STORE_ZJ_230_Split/split_req
      -- CP-element group 0: 	 assign_stmt_232/STORE_ZJ_230_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_232/STORE_ZJ_230_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_232/STORE_ZJ_230_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_232/STORE_ZJ_230_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_232/STORE_ZJ_230_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group initial_CP_1047_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:STORE_ZJ_230_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:STORE_ZJ_230_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    cr_1084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(0), ack => STORE_ZJ_230_store_0_req_1); -- 
    rr_1073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(0), ack => STORE_ZJ_230_store_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_232/STORE_ZJ_230_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_232/STORE_ZJ_230_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_232/STORE_ZJ_230_sample_completed_
      -- CP-element group 1: 	 assign_stmt_232/STORE_ZJ_230_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_232/STORE_ZJ_230_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initial_CP_1047_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:STORE_ZJ_230_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_ZJ_230_store_0_ack_0, ack => initial_CP_1047_elements(1)); -- 
    -- CP-element group 2:  branch  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	72 
    -- CP-element group 2:  members (13) 
      -- CP-element group 2: 	 assign_stmt_232/STORE_ZJ_230_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_233/branch_block_stmt_233__entry__
      -- CP-element group 2: 	 branch_block_stmt_233/merge_stmt_234__entry__
      -- CP-element group 2: 	 assign_stmt_232/STORE_ZJ_230_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_233/$entry
      -- CP-element group 2: 	 assign_stmt_232/$exit
      -- CP-element group 2: 	 assign_stmt_232/STORE_ZJ_230_Update/$exit
      -- CP-element group 2: 	 assign_stmt_232/STORE_ZJ_230_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_232/STORE_ZJ_230_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 branch_block_stmt_233/merge_stmt_234_dead_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_233/merge_stmt_234__entry___PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_233/merge_stmt_234__entry___PhiReq/phi_stmt_235/$entry
      -- CP-element group 2: 	 branch_block_stmt_233/merge_stmt_234__entry___PhiReq/phi_stmt_235/phi_stmt_235_sources/$entry
      -- 
    -- logger for CP element group initial_CP_1047_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:STORE_ZJ_230_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_ZJ_230_store_0_ack_1, ack => initial_CP_1047_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	77 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_233/assign_stmt_245/MUL_u12_u12_244_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_233/assign_stmt_245/MUL_u12_u12_244_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_233/assign_stmt_245/MUL_u12_u12_244_Sample/ra
      -- 
    -- logger for CP element group initial_CP_1047_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:MUL_u12_u12_244_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_u12_u12_244_inst_ack_0, ack => initial_CP_1047_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	77 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_233/assign_stmt_245/MUL_u12_u12_244_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_233/assign_stmt_245/MUL_u12_u12_244_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_233/assign_stmt_245/MUL_u12_u12_244_Update/ca
      -- 
    -- logger for CP element group initial_CP_1047_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:MUL_u12_u12_244_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_u12_u12_244_inst_ack_1, ack => initial_CP_1047_elements(4)); -- 
    -- CP-element group 5:  join  transition  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: 	77 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (9) 
      -- CP-element group 5: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_Sample/word_access_start/$entry
      -- CP-element group 5: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_Sample/word_access_start/word_0/rr
      -- CP-element group 5: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_Sample/word_access_start/word_0/$entry
      -- CP-element group 5: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_Sample/STORE_ZJ_241_Split/split_ack
      -- CP-element group 5: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_Sample/STORE_ZJ_241_Split/$exit
      -- CP-element group 5: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_Sample/STORE_ZJ_241_Split/split_req
      -- CP-element group 5: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_Sample/STORE_ZJ_241_Split/$entry
      -- CP-element group 5: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_sample_start_
      -- 
    -- logger for CP element group initial_CP_1047_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:STORE_ZJ_241_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(5), ack => STORE_ZJ_241_store_0_req_0); -- 
    initial_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "initial_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(4) & initial_CP_1047_elements(77);
      gj_initial_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (5) 
      -- CP-element group 6: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_Sample/word_access_start/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_Sample/word_access_start/word_0/ra
      -- CP-element group 6: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_Sample/word_access_start/$exit
      -- CP-element group 6: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_sample_completed_
      -- 
    -- logger for CP element group initial_CP_1047_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:STORE_ZJ_241_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_ZJ_241_store_0_ack_0, ack => initial_CP_1047_elements(6)); -- 
    -- CP-element group 7:  transition  place  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	77 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	9 
    -- CP-element group 7:  members (11) 
      -- CP-element group 7: 	 branch_block_stmt_233/assign_stmt_245__exit__
      -- CP-element group 7: 	 branch_block_stmt_233/branch_block_stmt_246__entry__
      -- CP-element group 7: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_Update/word_access_complete/$exit
      -- CP-element group 7: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_Update/word_access_complete/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_Update/word_access_complete/word_0/ca
      -- CP-element group 7: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_233/assign_stmt_245/$exit
      -- CP-element group 7: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247__entry__
      -- CP-element group 7: 	 branch_block_stmt_233/branch_block_stmt_246/branch_block_stmt_246__entry__
      -- CP-element group 7: 	 branch_block_stmt_233/branch_block_stmt_246/$entry
      -- CP-element group 7: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_Update/$exit
      -- 
    -- logger for CP element group initial_CP_1047_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:STORE_ZJ_241_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_ZJ_241_store_0_ack_1, ack => initial_CP_1047_elements(7)); -- 
    -- CP-element group 8:  fork  transition  place  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	67 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	68 
    -- CP-element group 8: 	69 
    -- CP-element group 8:  members (12) 
      -- CP-element group 8: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247__exit__
      -- CP-element group 8: 	 branch_block_stmt_233/branch_block_stmt_246__exit__
      -- CP-element group 8: 	 branch_block_stmt_233/assign_stmt_290__entry__
      -- CP-element group 8: 	 branch_block_stmt_233/branch_block_stmt_246/branch_block_stmt_246__exit__
      -- CP-element group 8: 	 branch_block_stmt_233/branch_block_stmt_246/$exit
      -- CP-element group 8: 	 branch_block_stmt_233/assign_stmt_290/$entry
      -- CP-element group 8: 	 branch_block_stmt_233/assign_stmt_290/ADD_u12_u12_289_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_233/assign_stmt_290/ADD_u12_u12_289_update_start_
      -- CP-element group 8: 	 branch_block_stmt_233/assign_stmt_290/ADD_u12_u12_289_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_233/assign_stmt_290/ADD_u12_u12_289_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_233/assign_stmt_290/ADD_u12_u12_289_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_233/assign_stmt_290/ADD_u12_u12_289_Update/cr
      -- 
    -- logger for CP element group initial_CP_1047_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:ADD_u12_u12_289_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:ADD_u12_u12_289_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    rr_1359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(8), ack => ADD_u12_u12_289_inst_req_0); -- 
    cr_1364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(8), ack => ADD_u12_u12_289_inst_req_1); -- 
    initial_CP_1047_elements(8) <= initial_CP_1047_elements(67);
    -- CP-element group 9:  transition  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	7 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	15 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247__entry__
      -- CP-element group 9: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/$entry
      -- 
    -- logger for CP element group initial_CP_1047_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    initial_CP_1047_elements(9) <= initial_CP_1047_elements(7);
    -- CP-element group 10:  merge  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	67 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247__exit__
      -- 
    -- logger for CP element group initial_CP_1047_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(10) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initial_CP_1047_elements(10) is bound as output of CP function.
    -- CP-element group 11:  merge  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/loop_back
      -- 
    -- logger for CP element group initial_CP_1047_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initial_CP_1047_elements(11) is bound as output of CP function.
    -- CP-element group 12:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	65 
    -- CP-element group 12: 	66 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/condition_done
      -- CP-element group 12: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/loop_exit/$entry
      -- CP-element group 12: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/loop_taken/$entry
      -- 
    -- logger for CP element group initial_CP_1047_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    initial_CP_1047_elements(12) <= initial_CP_1047_elements(17);
    -- CP-element group 13:  branch  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	59 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/loop_body_done
      -- 
    -- logger for CP element group initial_CP_1047_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    initial_CP_1047_elements(13) <= initial_CP_1047_elements(59);
    -- CP-element group 14:  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	23 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group initial_CP_1047_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    initial_CP_1047_elements(14) <= initial_CP_1047_elements(11);
    -- CP-element group 15:  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	25 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group initial_CP_1047_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(15) fired."); 
        -- 
      end if; --
    end process; 
    initial_CP_1047_elements(15) <= initial_CP_1047_elements(9);
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	19 
    -- CP-element group 16: 	20 
    -- CP-element group 16: 	46 
    -- CP-element group 16: 	64 
    -- CP-element group 16:  members (4) 
      -- CP-element group 16: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/loop_body_start
      -- CP-element group 16: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/$entry
      -- CP-element group 16: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_word_address_calculated
      -- CP-element group 16: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_root_address_calculated
      -- 
    -- logger for CP element group initial_CP_1047_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(16) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initial_CP_1047_elements(16) is bound as output of CP function.
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	22 
    -- CP-element group 17: 	63 
    -- CP-element group 17: 	64 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/condition_evaluated
      -- 
    -- logger for CP element group initial_CP_1047_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:do_while_stmt_247_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_1172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(17), ack => do_while_stmt_247_branch_req_0); -- 
    initial_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "initial_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initial_CP_1047_elements(22) & initial_CP_1047_elements(63) & initial_CP_1047_elements(64);
      gj_initial_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	22 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/aggregated_phi_sample_req
      -- CP-element group 18: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/phi_stmt_249_sample_start__ps
      -- 
    -- logger for CP element group initial_CP_1047_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(18) fired."); 
        -- 
      end if; --
    end process; 
    initial_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "initial_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(19) & initial_CP_1047_elements(22);
      gj_initial_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	16 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	21 
    -- CP-element group 19: 	63 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	18 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/phi_stmt_249_sample_start_
      -- 
    -- logger for CP element group initial_CP_1047_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(19) fired."); 
        -- 
      end if; --
    end process; 
    initial_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 27) := "initial_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initial_CP_1047_elements(16) & initial_CP_1047_elements(21) & initial_CP_1047_elements(63);
      gj_initial_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	16 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	22 
    -- CP-element group 20: 	38 
    -- CP-element group 20: 	42 
    -- CP-element group 20: 	62 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/aggregated_phi_update_req
      -- CP-element group 20: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/phi_stmt_249_update_start__ps
      -- CP-element group 20: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/phi_stmt_249_update_start_
      -- 
    -- logger for CP element group initial_CP_1047_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(20) fired."); 
        -- 
      end if; --
    end process; 
    initial_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "initial_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= initial_CP_1047_elements(16) & initial_CP_1047_elements(22) & initial_CP_1047_elements(38) & initial_CP_1047_elements(42) & initial_CP_1047_elements(62);
      gj_initial_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	61 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	19 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/phi_stmt_249_sample_completed__ps
      -- CP-element group 21: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/aggregated_phi_sample_ack
      -- CP-element group 21: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/phi_stmt_249_sample_completed_
      -- 
    -- logger for CP element group initial_CP_1047_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(21) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initial_CP_1047_elements(21) is bound as output of CP function.
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	17 
    -- CP-element group 22: 	36 
    -- CP-element group 22: 	40 
    -- CP-element group 22: 	60 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	18 
    -- CP-element group 22: 	20 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/phi_stmt_249_update_completed__ps
      -- CP-element group 22: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/phi_stmt_249_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/aggregated_phi_update_ack
      -- 
    -- logger for CP element group initial_CP_1047_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(22) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initial_CP_1047_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	14 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/phi_stmt_249_loopback_trigger
      -- 
    -- logger for CP element group initial_CP_1047_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(23) fired."); 
        -- 
      end if; --
    end process; 
    initial_CP_1047_elements(23) <= initial_CP_1047_elements(14);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/phi_stmt_249_loopback_sample_req
      -- CP-element group 24: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/phi_stmt_249_loopback_sample_req_ps
      -- 
    -- logger for CP element group initial_CP_1047_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:phi_stmt_249_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_249_loopback_sample_req_1187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_249_loopback_sample_req_1187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(24), ack => phi_stmt_249_req_1); -- 
    -- Element group initial_CP_1047_elements(24) is bound as output of CP function.
    -- CP-element group 25:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	15 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/phi_stmt_249_entry_trigger
      -- 
    -- logger for CP element group initial_CP_1047_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(25) fired."); 
        -- 
      end if; --
    end process; 
    initial_CP_1047_elements(25) <= initial_CP_1047_elements(15);
    -- CP-element group 26:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/phi_stmt_249_entry_sample_req
      -- CP-element group 26: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/phi_stmt_249_entry_sample_req_ps
      -- 
    -- logger for CP element group initial_CP_1047_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:phi_stmt_249_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_249_entry_sample_req_1190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_249_entry_sample_req_1190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(26), ack => phi_stmt_249_req_0); -- 
    -- Element group initial_CP_1047_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/phi_stmt_249_phi_mux_ack_ps
      -- CP-element group 27: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/phi_stmt_249_phi_mux_ack
      -- 
    -- logger for CP element group initial_CP_1047_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:phi_stmt_249_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_249_phi_mux_ack_1193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_249_ack_0, ack => initial_CP_1047_elements(27)); -- 
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_252_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_252_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_252_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_252_sample_completed_
      -- 
    -- logger for CP element group initial_CP_1047_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(28) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initial_CP_1047_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_252_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_252_update_start_
      -- 
    -- logger for CP element group initial_CP_1047_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(29) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initial_CP_1047_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_252_update_completed__ps
      -- 
    -- logger for CP element group initial_CP_1047_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(30) fired."); 
        -- 
      end if; --
    end process; 
    initial_CP_1047_elements(30) <= initial_CP_1047_elements(31);
    -- CP-element group 31:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	30 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_252_update_completed_
      -- 
    -- logger for CP element group initial_CP_1047_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(31) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initial_CP_1047_elements(31) is a control-delay.
    cp_element_31_delay: control_delay_element  generic map(name => " 31_delay", delay_value => 1)  port map(req => initial_CP_1047_elements(29), ack => initial_CP_1047_elements(31), clk => clk, reset =>reset);
    -- CP-element group 32:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/R_NI_253_Sample/req
      -- CP-element group 32: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/R_NI_253_sample_start__ps
      -- CP-element group 32: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/R_NI_253_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/R_NI_253_Sample/$entry
      -- 
    -- logger for CP element group initial_CP_1047_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:NI_280_253_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(32), ack => NI_280_253_buf_req_0); -- 
    -- Element group initial_CP_1047_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/R_NI_253_update_start__ps
      -- CP-element group 33: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/R_NI_253_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/R_NI_253_Update/req
      -- CP-element group 33: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/R_NI_253_update_start_
      -- 
    -- logger for CP element group initial_CP_1047_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:NI_280_253_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(33), ack => NI_280_253_buf_req_1); -- 
    -- Element group initial_CP_1047_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/R_NI_253_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/R_NI_253_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/R_NI_253_Sample/ack
      -- CP-element group 34: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/R_NI_253_sample_completed__ps
      -- 
    -- logger for CP element group initial_CP_1047_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:NI_280_253_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NI_280_253_buf_ack_0, ack => initial_CP_1047_elements(34)); -- 
    -- CP-element group 35:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/R_NI_253_update_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/R_NI_253_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/R_NI_253_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/R_NI_253_Update/ack
      -- 
    -- logger for CP element group initial_CP_1047_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:NI_280_253_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NI_280_253_buf_ack_1, ack => initial_CP_1047_elements(35)); -- 
    -- CP-element group 36:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	22 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	38 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_257_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_257_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_257_Sample/rr
      -- 
    -- logger for CP element group initial_CP_1047_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(36) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:type_cast_257_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(36), ack => type_cast_257_inst_req_0); -- 
    initial_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "initial_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(22) & initial_CP_1047_elements(38);
      gj_initial_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: 	54 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_257_update_start_
      -- CP-element group 37: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_257_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_257_Update/cr
      -- 
    -- logger for CP element group initial_CP_1047_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:type_cast_257_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(37), ack => type_cast_257_inst_req_1); -- 
    initial_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "initial_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(39) & initial_CP_1047_elements(54);
      gj_initial_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	20 
    -- CP-element group 38: 	36 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_257_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_257_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_257_Sample/ra
      -- 
    -- logger for CP element group initial_CP_1047_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(38) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:type_cast_257_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_257_inst_ack_0, ack => initial_CP_1047_elements(38)); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	52 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_257_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_257_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_257_Update/ca
      -- 
    -- logger for CP element group initial_CP_1047_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:type_cast_257_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_257_inst_ack_1, ack => initial_CP_1047_elements(39)); -- 
    -- CP-element group 40:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	22 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	42 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_261_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_261_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_261_Sample/req
      -- 
    -- logger for CP element group initial_CP_1047_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(40) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:W_I_230_delayed_4_0_259_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(40), ack => W_I_230_delayed_4_0_259_inst_req_0); -- 
    initial_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "initial_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(22) & initial_CP_1047_elements(42);
      gj_initial_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	43 
    -- CP-element group 41: 	50 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_261_update_start_
      -- CP-element group 41: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_261_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_261_Update/req
      -- 
    -- logger for CP element group initial_CP_1047_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(41) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:W_I_230_delayed_4_0_259_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(41), ack => W_I_230_delayed_4_0_259_inst_req_1); -- 
    initial_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "initial_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(43) & initial_CP_1047_elements(50);
      gj_initial_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: marked-successors 
    -- CP-element group 42: 	20 
    -- CP-element group 42: 	40 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_261_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_261_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_261_Sample/ack
      -- 
    -- logger for CP element group initial_CP_1047_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(42) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:W_I_230_delayed_4_0_259_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_I_230_delayed_4_0_259_inst_ack_0, ack => initial_CP_1047_elements(42)); -- 
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	41 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_261_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_261_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_261_Update/ack
      -- 
    -- logger for CP element group initial_CP_1047_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(43) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:W_I_230_delayed_4_0_259_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_I_230_delayed_4_0_259_inst_ack_1, ack => initial_CP_1047_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: 	49 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	50 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	50 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_266_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_266_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_266_Sample/rr
      -- 
    -- logger for CP element group initial_CP_1047_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(44) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:type_cast_266_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(44), ack => type_cast_266_inst_req_0); -- 
    initial_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "initial_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initial_CP_1047_elements(43) & initial_CP_1047_elements(49) & initial_CP_1047_elements(50);
      gj_initial_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: marked-predecessors 
    -- CP-element group 45: 	51 
    -- CP-element group 45: 	58 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	51 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_266_update_start_
      -- CP-element group 45: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_266_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_266_Update/cr
      -- 
    -- logger for CP element group initial_CP_1047_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(45) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:type_cast_266_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(45), ack => type_cast_266_inst_req_1); -- 
    initial_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "initial_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(51) & initial_CP_1047_elements(58);
      gj_initial_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	16 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	48 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (5) 
      -- CP-element group 46: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_Sample/word_access_start/$entry
      -- CP-element group 46: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_Sample/word_access_start/word_0/$entry
      -- CP-element group 46: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initial_CP_1047_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(46) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:LOAD_ZJ_263_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(46), ack => LOAD_ZJ_263_load_0_req_0); -- 
    initial_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "initial_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(16) & initial_CP_1047_elements(48);
      gj_initial_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	49 
    -- CP-element group 47: 	50 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (5) 
      -- CP-element group 47: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_update_start_
      -- CP-element group 47: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_Update/$entry
      -- CP-element group 47: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_Update/word_access_complete/$entry
      -- CP-element group 47: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_Update/word_access_complete/word_0/$entry
      -- CP-element group 47: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group initial_CP_1047_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(47) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:LOAD_ZJ_263_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(47), ack => LOAD_ZJ_263_load_0_req_1); -- 
    initial_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "initial_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(49) & initial_CP_1047_elements(50);
      gj_initial_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: marked-successors 
    -- CP-element group 48: 	46 
    -- CP-element group 48:  members (5) 
      -- CP-element group 48: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_Sample/word_access_start/$exit
      -- CP-element group 48: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_Sample/word_access_start/word_0/$exit
      -- CP-element group 48: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initial_CP_1047_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(48) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:LOAD_ZJ_263_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ZJ_263_load_0_ack_0, ack => initial_CP_1047_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	44 
    -- CP-element group 49: marked-successors 
    -- CP-element group 49: 	47 
    -- CP-element group 49:  members (9) 
      -- CP-element group 49: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_Update/word_access_complete/$exit
      -- CP-element group 49: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_Update/word_access_complete/word_0/$exit
      -- CP-element group 49: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_Update/word_access_complete/word_0/ca
      -- CP-element group 49: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_Update/LOAD_ZJ_263_Merge/$entry
      -- CP-element group 49: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_Update/LOAD_ZJ_263_Merge/$exit
      -- CP-element group 49: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_Update/LOAD_ZJ_263_Merge/merge_req
      -- CP-element group 49: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/LOAD_ZJ_263_Update/LOAD_ZJ_263_Merge/merge_ack
      -- 
    -- logger for CP element group initial_CP_1047_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(49) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:LOAD_ZJ_263_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ZJ_263_load_0_ack_1, ack => initial_CP_1047_elements(49)); -- 
    -- CP-element group 50:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	44 
    -- CP-element group 50: successors 
    -- CP-element group 50: marked-successors 
    -- CP-element group 50: 	41 
    -- CP-element group 50: 	44 
    -- CP-element group 50: 	47 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_266_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_266_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_266_Sample/ra
      -- 
    -- logger for CP element group initial_CP_1047_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(50) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:type_cast_266_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_266_inst_ack_0, ack => initial_CP_1047_elements(50)); -- 
    -- CP-element group 51:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	45 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	56 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	45 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_266_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_266_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/type_cast_266_Update/ca
      -- 
    -- logger for CP element group initial_CP_1047_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(51) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:type_cast_266_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_266_inst_ack_1, ack => initial_CP_1047_elements(51)); -- 
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	39 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_270_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_270_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_270_Sample/req
      -- 
    -- logger for CP element group initial_CP_1047_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(52) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:W_wdata_236_delayed_4_0_268_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(52), ack => W_wdata_236_delayed_4_0_268_inst_req_0); -- 
    initial_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "initial_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(39) & initial_CP_1047_elements(54);
      gj_initial_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	55 
    -- CP-element group 53: 	58 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_270_update_start_
      -- CP-element group 53: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_270_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_270_Update/req
      -- 
    -- logger for CP element group initial_CP_1047_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(53) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:W_wdata_236_delayed_4_0_268_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(53), ack => W_wdata_236_delayed_4_0_268_inst_req_1); -- 
    initial_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "initial_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(55) & initial_CP_1047_elements(58);
      gj_initial_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	37 
    -- CP-element group 54: 	52 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_270_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_270_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_270_Sample/ack
      -- 
    -- logger for CP element group initial_CP_1047_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(54) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:W_wdata_236_delayed_4_0_268_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_236_delayed_4_0_268_inst_ack_0, ack => initial_CP_1047_elements(54)); -- 
    -- CP-element group 55:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: marked-successors 
    -- CP-element group 55: 	53 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_270_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_270_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/assign_stmt_270_Update/ack
      -- 
    -- logger for CP element group initial_CP_1047_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(55) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:W_wdata_236_delayed_4_0_268_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_236_delayed_4_0_268_inst_ack_1, ack => initial_CP_1047_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	51 
    -- CP-element group 56: 	55 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/call_stmt_275_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/call_stmt_275_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/call_stmt_275_Sample/crr
      -- 
    -- logger for CP element group initial_CP_1047_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(56) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:call_stmt_275_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(56), ack => call_stmt_275_call_req_0); -- 
    initial_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "initial_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initial_CP_1047_elements(51) & initial_CP_1047_elements(55) & initial_CP_1047_elements(58);
      gj_initial_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	59 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/call_stmt_275_update_start_
      -- CP-element group 57: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/call_stmt_275_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/call_stmt_275_Update/ccr
      -- 
    -- logger for CP element group initial_CP_1047_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(57) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:call_stmt_275_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_1323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(57), ack => call_stmt_275_call_req_1); -- 
    initial_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "initial_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= initial_CP_1047_elements(59);
      gj_initial_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	53 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/call_stmt_275_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/call_stmt_275_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/call_stmt_275_Sample/cra
      -- 
    -- logger for CP element group initial_CP_1047_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(58) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:call_stmt_275_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_275_call_ack_0, ack => initial_CP_1047_elements(58)); -- 
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	13 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	57 
    -- CP-element group 59:  members (4) 
      -- CP-element group 59: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/$exit
      -- CP-element group 59: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/call_stmt_275_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/call_stmt_275_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/call_stmt_275_Update/cca
      -- 
    -- logger for CP element group initial_CP_1047_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(59) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:call_stmt_275_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_275_call_ack_1, ack => initial_CP_1047_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	22 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/ADD_u12_u12_279_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/ADD_u12_u12_279_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/ADD_u12_u12_279_Sample/rr
      -- 
    -- logger for CP element group initial_CP_1047_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(60) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:ADD_u12_u12_279_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(60), ack => ADD_u12_u12_279_inst_req_0); -- 
    initial_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "initial_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(22) & initial_CP_1047_elements(62);
      gj_initial_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	21 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/ADD_u12_u12_279_update_start_
      -- CP-element group 61: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/ADD_u12_u12_279_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/ADD_u12_u12_279_Update/cr
      -- 
    -- logger for CP element group initial_CP_1047_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(61) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:ADD_u12_u12_279_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(61), ack => ADD_u12_u12_279_inst_req_1); -- 
    initial_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "initial_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(21) & initial_CP_1047_elements(63);
      gj_initial_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	20 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/ADD_u12_u12_279_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/ADD_u12_u12_279_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/ADD_u12_u12_279_Sample/ra
      -- 
    -- logger for CP element group initial_CP_1047_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(62) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:ADD_u12_u12_279_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_279_inst_ack_0, ack => initial_CP_1047_elements(62)); -- 
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	17 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	19 
    -- CP-element group 63: 	61 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/ADD_u12_u12_279_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/ADD_u12_u12_279_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/ADD_u12_u12_279_Update/ca
      -- 
    -- logger for CP element group initial_CP_1047_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(63) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:ADD_u12_u12_279_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_279_inst_ack_1, ack => initial_CP_1047_elements(63)); -- 
    -- CP-element group 64:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	16 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	17 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/do_while_stmt_247_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group initial_CP_1047_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(64) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initial_CP_1047_elements(64) is a control-delay.
    cp_element_64_delay: control_delay_element  generic map(name => " 64_delay", delay_value => 1)  port map(req => initial_CP_1047_elements(16), ack => initial_CP_1047_elements(64), clk => clk, reset =>reset);
    -- CP-element group 65:  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	12 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/loop_exit/$exit
      -- CP-element group 65: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/loop_exit/ack
      -- 
    -- logger for CP element group initial_CP_1047_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(65) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:do_while_stmt_247_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_247_branch_ack_0, ack => initial_CP_1047_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	12 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/loop_taken/$exit
      -- CP-element group 66: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/loop_taken/ack
      -- 
    -- logger for CP element group initial_CP_1047_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(66) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:do_while_stmt_247_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_247_branch_ack_1, ack => initial_CP_1047_elements(66)); -- 
    -- CP-element group 67:  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	10 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	8 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_233/branch_block_stmt_246/do_while_stmt_247/$exit
      -- 
    -- logger for CP element group initial_CP_1047_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(67) fired."); 
        -- 
      end if; --
    end process; 
    initial_CP_1047_elements(67) <= initial_CP_1047_elements(10);
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	8 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_233/assign_stmt_290/ADD_u12_u12_289_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_233/assign_stmt_290/ADD_u12_u12_289_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_233/assign_stmt_290/ADD_u12_u12_289_Sample/ra
      -- 
    -- logger for CP element group initial_CP_1047_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(68) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:ADD_u12_u12_289_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_289_inst_ack_0, ack => initial_CP_1047_elements(68)); -- 
    -- CP-element group 69:  branch  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	8 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (27) 
      -- CP-element group 69: 	 branch_block_stmt_233/assign_stmt_290__exit__
      -- CP-element group 69: 	 branch_block_stmt_233/if_stmt_291__entry__
      -- CP-element group 69: 	 branch_block_stmt_233/assign_stmt_290/$exit
      -- CP-element group 69: 	 branch_block_stmt_233/assign_stmt_290/ADD_u12_u12_289_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_233/assign_stmt_290/ADD_u12_u12_289_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_233/assign_stmt_290/ADD_u12_u12_289_Update/ca
      -- CP-element group 69: 	 branch_block_stmt_233/if_stmt_291_dead_link/$entry
      -- CP-element group 69: 	 branch_block_stmt_233/if_stmt_291_eval_test/$entry
      -- CP-element group 69: 	 branch_block_stmt_233/if_stmt_291_eval_test/$exit
      -- CP-element group 69: 	 branch_block_stmt_233/if_stmt_291_eval_test/ULT_u12_u1_294/$entry
      -- CP-element group 69: 	 branch_block_stmt_233/if_stmt_291_eval_test/ULT_u12_u1_294/$exit
      -- CP-element group 69: 	 branch_block_stmt_233/if_stmt_291_eval_test/ULT_u12_u1_294/ULT_u12_u1_294_inputs/$entry
      -- CP-element group 69: 	 branch_block_stmt_233/if_stmt_291_eval_test/ULT_u12_u1_294/ULT_u12_u1_294_inputs/$exit
      -- CP-element group 69: 	 branch_block_stmt_233/if_stmt_291_eval_test/ULT_u12_u1_294/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_233/if_stmt_291_eval_test/ULT_u12_u1_294/SplitProtocol/$exit
      -- CP-element group 69: 	 branch_block_stmt_233/if_stmt_291_eval_test/ULT_u12_u1_294/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_233/if_stmt_291_eval_test/ULT_u12_u1_294/SplitProtocol/Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_233/if_stmt_291_eval_test/ULT_u12_u1_294/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_233/if_stmt_291_eval_test/ULT_u12_u1_294/SplitProtocol/Sample/ra
      -- CP-element group 69: 	 branch_block_stmt_233/if_stmt_291_eval_test/ULT_u12_u1_294/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_233/if_stmt_291_eval_test/ULT_u12_u1_294/SplitProtocol/Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_233/if_stmt_291_eval_test/ULT_u12_u1_294/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_233/if_stmt_291_eval_test/ULT_u12_u1_294/SplitProtocol/Update/ca
      -- CP-element group 69: 	 branch_block_stmt_233/if_stmt_291_eval_test/branch_req
      -- CP-element group 69: 	 branch_block_stmt_233/ULT_u12_u1_294_place
      -- CP-element group 69: 	 branch_block_stmt_233/if_stmt_291_if_link/$entry
      -- CP-element group 69: 	 branch_block_stmt_233/if_stmt_291_else_link/$entry
      -- 
    -- logger for CP element group initial_CP_1047_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(69) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:ADD_u12_u12_289_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:if_stmt_291_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_1365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_289_inst_ack_1, ack => initial_CP_1047_elements(69)); -- 
    branch_req_1392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(69), ack => if_stmt_291_branch_req_0); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	73 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (11) 
      -- CP-element group 70: 	 branch_block_stmt_233/if_stmt_291_if_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_233/if_stmt_291_if_link/if_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_233/loopback
      -- CP-element group 70: 	 branch_block_stmt_233/loopback_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_233/loopback_PhiReq/phi_stmt_235/$entry
      -- CP-element group 70: 	 branch_block_stmt_233/loopback_PhiReq/phi_stmt_235/phi_stmt_235_sources/$entry
      -- CP-element group 70: 	 branch_block_stmt_233/loopback_PhiReq/phi_stmt_235/phi_stmt_235_sources/Interlock/$entry
      -- CP-element group 70: 	 branch_block_stmt_233/loopback_PhiReq/phi_stmt_235/phi_stmt_235_sources/Interlock/Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_233/loopback_PhiReq/phi_stmt_235/phi_stmt_235_sources/Interlock/Sample/req
      -- CP-element group 70: 	 branch_block_stmt_233/loopback_PhiReq/phi_stmt_235/phi_stmt_235_sources/Interlock/Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_233/loopback_PhiReq/phi_stmt_235/phi_stmt_235_sources/Interlock/Update/req
      -- 
    -- logger for CP element group initial_CP_1047_elements(70)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(70)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(70) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:if_stmt_291_branch_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:YI_290_239_buf_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:YI_290_239_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_1397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_291_branch_ack_1, ack => initial_CP_1047_elements(70)); -- 
    req_1433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(70), ack => YI_290_239_buf_req_0); -- 
    req_1438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(70), ack => YI_290_239_buf_req_1); -- 
    -- CP-element group 71:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	78 
    -- CP-element group 71: 	79 
    -- CP-element group 71:  members (22) 
      -- CP-element group 71: 	 branch_block_stmt_233/branch_block_stmt_233__exit__
      -- CP-element group 71: 	 branch_block_stmt_233/$exit
      -- CP-element group 71: 	 branch_block_stmt_233/if_stmt_291__exit__
      -- CP-element group 71: 	 branch_block_stmt_233/if_stmt_291_else_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_233/if_stmt_291_else_link/else_choice_transition
      -- CP-element group 71: 	 assign_stmt_300/$entry
      -- CP-element group 71: 	 assign_stmt_300/STORE_ZJ_298_sample_start_
      -- CP-element group 71: 	 assign_stmt_300/STORE_ZJ_298_update_start_
      -- CP-element group 71: 	 assign_stmt_300/STORE_ZJ_298_word_address_calculated
      -- CP-element group 71: 	 assign_stmt_300/STORE_ZJ_298_root_address_calculated
      -- CP-element group 71: 	 assign_stmt_300/STORE_ZJ_298_Sample/$entry
      -- CP-element group 71: 	 assign_stmt_300/STORE_ZJ_298_Sample/STORE_ZJ_298_Split/$entry
      -- CP-element group 71: 	 assign_stmt_300/STORE_ZJ_298_Sample/STORE_ZJ_298_Split/$exit
      -- CP-element group 71: 	 assign_stmt_300/STORE_ZJ_298_Sample/STORE_ZJ_298_Split/split_req
      -- CP-element group 71: 	 assign_stmt_300/STORE_ZJ_298_Sample/STORE_ZJ_298_Split/split_ack
      -- CP-element group 71: 	 assign_stmt_300/STORE_ZJ_298_Sample/word_access_start/$entry
      -- CP-element group 71: 	 assign_stmt_300/STORE_ZJ_298_Sample/word_access_start/word_0/$entry
      -- CP-element group 71: 	 assign_stmt_300/STORE_ZJ_298_Sample/word_access_start/word_0/rr
      -- CP-element group 71: 	 assign_stmt_300/STORE_ZJ_298_Update/$entry
      -- CP-element group 71: 	 assign_stmt_300/STORE_ZJ_298_Update/word_access_complete/$entry
      -- CP-element group 71: 	 assign_stmt_300/STORE_ZJ_298_Update/word_access_complete/word_0/$entry
      -- CP-element group 71: 	 assign_stmt_300/STORE_ZJ_298_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group initial_CP_1047_elements(71)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(71)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(71) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:if_stmt_291_branch_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:STORE_ZJ_298_store_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:STORE_ZJ_298_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_1401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_291_branch_ack_0, ack => initial_CP_1047_elements(71)); -- 
    rr_1469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(71), ack => STORE_ZJ_298_store_0_req_0); -- 
    cr_1480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(71), ack => STORE_ZJ_298_store_0_req_1); -- 
    -- CP-element group 72:  transition  output  delay-element  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	2 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	76 
    -- CP-element group 72:  members (5) 
      -- CP-element group 72: 	 branch_block_stmt_233/merge_stmt_234__entry___PhiReq/$exit
      -- CP-element group 72: 	 branch_block_stmt_233/merge_stmt_234__entry___PhiReq/phi_stmt_235/$exit
      -- CP-element group 72: 	 branch_block_stmt_233/merge_stmt_234__entry___PhiReq/phi_stmt_235/phi_stmt_235_sources/$exit
      -- CP-element group 72: 	 branch_block_stmt_233/merge_stmt_234__entry___PhiReq/phi_stmt_235/phi_stmt_235_sources/type_cast_238_konst_delay_trans
      -- CP-element group 72: 	 branch_block_stmt_233/merge_stmt_234__entry___PhiReq/phi_stmt_235/phi_stmt_235_req
      -- 
    -- logger for CP element group initial_CP_1047_elements(72)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(72)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(72) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:phi_stmt_235_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_235_req_1417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_235_req_1417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(72), ack => phi_stmt_235_req_0); -- 
    -- Element group initial_CP_1047_elements(72) is a control-delay.
    cp_element_72_delay: control_delay_element  generic map(name => " 72_delay", delay_value => 1)  port map(req => initial_CP_1047_elements(2), ack => initial_CP_1047_elements(72), clk => clk, reset =>reset);
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	70 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_233/loopback_PhiReq/phi_stmt_235/phi_stmt_235_sources/Interlock/Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_233/loopback_PhiReq/phi_stmt_235/phi_stmt_235_sources/Interlock/Sample/ack
      -- 
    -- logger for CP element group initial_CP_1047_elements(73)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(73)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(73) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:YI_290_239_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => YI_290_239_buf_ack_0, ack => initial_CP_1047_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_233/loopback_PhiReq/phi_stmt_235/phi_stmt_235_sources/Interlock/Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_233/loopback_PhiReq/phi_stmt_235/phi_stmt_235_sources/Interlock/Update/ack
      -- 
    -- logger for CP element group initial_CP_1047_elements(74)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(74)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(74) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:YI_290_239_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => YI_290_239_buf_ack_1, ack => initial_CP_1047_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_233/loopback_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_233/loopback_PhiReq/phi_stmt_235/$exit
      -- CP-element group 75: 	 branch_block_stmt_233/loopback_PhiReq/phi_stmt_235/phi_stmt_235_sources/$exit
      -- CP-element group 75: 	 branch_block_stmt_233/loopback_PhiReq/phi_stmt_235/phi_stmt_235_sources/Interlock/$exit
      -- CP-element group 75: 	 branch_block_stmt_233/loopback_PhiReq/phi_stmt_235/phi_stmt_235_req
      -- 
    -- logger for CP element group initial_CP_1047_elements(75)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(75)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(75) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:phi_stmt_235_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_235_req_1440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_235_req_1440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(75), ack => phi_stmt_235_req_1); -- 
    initial_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "initial_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(73) & initial_CP_1047_elements(74);
      gj_initial_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  merge  transition  place  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	72 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_233/merge_stmt_234_PhiReqMerge
      -- CP-element group 76: 	 branch_block_stmt_233/merge_stmt_234_PhiAck/$entry
      -- 
    -- logger for CP element group initial_CP_1047_elements(76)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(76)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(76) fired."); 
        -- 
      end if; --
    end process; 
    initial_CP_1047_elements(76) <= OrReduce(initial_CP_1047_elements(72) & initial_CP_1047_elements(75));
    -- CP-element group 77:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	3 
    -- CP-element group 77: 	4 
    -- CP-element group 77: 	5 
    -- CP-element group 77: 	7 
    -- CP-element group 77:  members (18) 
      -- CP-element group 77: 	 branch_block_stmt_233/merge_stmt_234__exit__
      -- CP-element group 77: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_update_start_
      -- CP-element group 77: 	 branch_block_stmt_233/assign_stmt_245__entry__
      -- CP-element group 77: 	 branch_block_stmt_233/assign_stmt_245/MUL_u12_u12_244_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_233/assign_stmt_245/MUL_u12_u12_244_update_start_
      -- CP-element group 77: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_233/assign_stmt_245/$entry
      -- CP-element group 77: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_233/assign_stmt_245/MUL_u12_u12_244_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_233/assign_stmt_245/MUL_u12_u12_244_Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_233/assign_stmt_245/MUL_u12_u12_244_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_233/assign_stmt_245/MUL_u12_u12_244_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_233/assign_stmt_245/STORE_ZJ_241_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_233/merge_stmt_234_PhiAck/$exit
      -- CP-element group 77: 	 branch_block_stmt_233/merge_stmt_234_PhiAck/phi_stmt_235_ack
      -- 
    -- logger for CP element group initial_CP_1047_elements(77)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(77)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(77) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:phi_stmt_235_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:STORE_ZJ_241_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:MUL_u12_u12_244_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:MUL_u12_u12_244_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_235_ack_1445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_235_ack_0, ack => initial_CP_1047_elements(77)); -- 
    cr_1149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(77), ack => STORE_ZJ_241_store_0_req_1); -- 
    rr_1111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(77), ack => MUL_u12_u12_244_inst_req_0); -- 
    cr_1116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(77), ack => MUL_u12_u12_244_inst_req_1); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	71 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 assign_stmt_300/STORE_ZJ_298_sample_completed_
      -- CP-element group 78: 	 assign_stmt_300/STORE_ZJ_298_Sample/$exit
      -- CP-element group 78: 	 assign_stmt_300/STORE_ZJ_298_Sample/word_access_start/$exit
      -- CP-element group 78: 	 assign_stmt_300/STORE_ZJ_298_Sample/word_access_start/word_0/$exit
      -- CP-element group 78: 	 assign_stmt_300/STORE_ZJ_298_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initial_CP_1047_elements(78)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(78)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(78) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:STORE_ZJ_298_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_ZJ_298_store_0_ack_0, ack => initial_CP_1047_elements(78)); -- 
    -- CP-element group 79:  transition  place  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	71 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (9) 
      -- CP-element group 79: 	 assign_stmt_300/$exit
      -- CP-element group 79: 	 assign_stmt_300/STORE_ZJ_298_update_completed_
      -- CP-element group 79: 	 assign_stmt_300/STORE_ZJ_298_Update/$exit
      -- CP-element group 79: 	 assign_stmt_300/STORE_ZJ_298_Update/word_access_complete/$exit
      -- CP-element group 79: 	 assign_stmt_300/STORE_ZJ_298_Update/word_access_complete/word_0/$exit
      -- CP-element group 79: 	 assign_stmt_300/STORE_ZJ_298_Update/word_access_complete/word_0/ca
      -- CP-element group 79: 	 branch_block_stmt_301/$entry
      -- CP-element group 79: 	 branch_block_stmt_301/branch_block_stmt_301__entry__
      -- CP-element group 79: 	 branch_block_stmt_301/do_while_stmt_302__entry__
      -- 
    -- logger for CP element group initial_CP_1047_elements(79)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(79)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(79) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:STORE_ZJ_298_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_ZJ_298_store_0_ack_1, ack => initial_CP_1047_elements(79)); -- 
    -- CP-element group 80:  transition  place  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	139 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 $exit
      -- CP-element group 80: 	 branch_block_stmt_301/$exit
      -- CP-element group 80: 	 branch_block_stmt_301/branch_block_stmt_301__exit__
      -- CP-element group 80: 	 branch_block_stmt_301/do_while_stmt_302__exit__
      -- 
    -- logger for CP element group initial_CP_1047_elements(80)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(80)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(80) fired."); 
        -- 
      end if; --
    end process; 
    initial_CP_1047_elements(80) <= initial_CP_1047_elements(139);
    -- CP-element group 81:  transition  place  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	87 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_301/do_while_stmt_302/$entry
      -- CP-element group 81: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302__entry__
      -- 
    -- logger for CP element group initial_CP_1047_elements(81)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(81)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(81) fired."); 
        -- 
      end if; --
    end process; 
    initial_CP_1047_elements(81) <= initial_CP_1047_elements(79);
    -- CP-element group 82:  merge  place  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	139 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302__exit__
      -- 
    -- logger for CP element group initial_CP_1047_elements(82)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(82)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(82) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initial_CP_1047_elements(82) is bound as output of CP function.
    -- CP-element group 83:  merge  place  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	86 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_301/do_while_stmt_302/loop_back
      -- 
    -- logger for CP element group initial_CP_1047_elements(83)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(83)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(83) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initial_CP_1047_elements(83) is bound as output of CP function.
    -- CP-element group 84:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	89 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	137 
    -- CP-element group 84: 	138 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_301/do_while_stmt_302/loop_taken/$entry
      -- CP-element group 84: 	 branch_block_stmt_301/do_while_stmt_302/condition_done
      -- CP-element group 84: 	 branch_block_stmt_301/do_while_stmt_302/loop_exit/$entry
      -- 
    -- logger for CP element group initial_CP_1047_elements(84)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(84)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(84) fired."); 
        -- 
      end if; --
    end process; 
    initial_CP_1047_elements(84) <= initial_CP_1047_elements(89);
    -- CP-element group 85:  branch  place  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	131 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_301/do_while_stmt_302/loop_body_done
      -- 
    -- logger for CP element group initial_CP_1047_elements(85)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(85)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(85) fired."); 
        -- 
      end if; --
    end process; 
    initial_CP_1047_elements(85) <= initial_CP_1047_elements(131);
    -- CP-element group 86:  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	83 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	95 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group initial_CP_1047_elements(86)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(86)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(86) fired."); 
        -- 
      end if; --
    end process; 
    initial_CP_1047_elements(86) <= initial_CP_1047_elements(83);
    -- CP-element group 87:  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	81 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	97 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group initial_CP_1047_elements(87)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(87)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(87) fired."); 
        -- 
      end if; --
    end process; 
    initial_CP_1047_elements(87) <= initial_CP_1047_elements(81);
    -- CP-element group 88:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	91 
    -- CP-element group 88: 	92 
    -- CP-element group 88: 	118 
    -- CP-element group 88: 	136 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/$entry
      -- CP-element group 88: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/loop_body_start
      -- CP-element group 88: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_word_address_calculated
      -- CP-element group 88: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_root_address_calculated
      -- 
    -- logger for CP element group initial_CP_1047_elements(88)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(88)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(88) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initial_CP_1047_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	94 
    -- CP-element group 89: 	135 
    -- CP-element group 89: 	136 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	84 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/condition_evaluated
      -- 
    -- logger for CP element group initial_CP_1047_elements(89)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(89)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(89) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:do_while_stmt_302_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_1503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(89), ack => do_while_stmt_302_branch_req_0); -- 
    initial_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "initial_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initial_CP_1047_elements(94) & initial_CP_1047_elements(135) & initial_CP_1047_elements(136);
      gj_initial_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	91 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	94 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/aggregated_phi_sample_req
      -- CP-element group 90: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/phi_stmt_304_sample_start__ps
      -- 
    -- logger for CP element group initial_CP_1047_elements(90)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(90)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(90) fired."); 
        -- 
      end if; --
    end process; 
    initial_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "initial_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(91) & initial_CP_1047_elements(94);
      gj_initial_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  join  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	88 
    -- CP-element group 91: marked-predecessors 
    -- CP-element group 91: 	93 
    -- CP-element group 91: 	135 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	90 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/phi_stmt_304_sample_start_
      -- 
    -- logger for CP element group initial_CP_1047_elements(91)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(91)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(91) fired."); 
        -- 
      end if; --
    end process; 
    initial_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 27) := "initial_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initial_CP_1047_elements(88) & initial_CP_1047_elements(93) & initial_CP_1047_elements(135);
      gj_initial_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	88 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	94 
    -- CP-element group 92: 	110 
    -- CP-element group 92: 	114 
    -- CP-element group 92: 	134 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/aggregated_phi_update_req
      -- CP-element group 92: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/phi_stmt_304_update_start_
      -- CP-element group 92: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/phi_stmt_304_update_start__ps
      -- 
    -- logger for CP element group initial_CP_1047_elements(92)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(92)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(92) fired."); 
        -- 
      end if; --
    end process; 
    initial_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "initial_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= initial_CP_1047_elements(88) & initial_CP_1047_elements(94) & initial_CP_1047_elements(110) & initial_CP_1047_elements(114) & initial_CP_1047_elements(134);
      gj_initial_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	133 
    -- CP-element group 93: marked-successors 
    -- CP-element group 93: 	91 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/aggregated_phi_sample_ack
      -- CP-element group 93: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/phi_stmt_304_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/phi_stmt_304_sample_completed__ps
      -- 
    -- logger for CP element group initial_CP_1047_elements(93)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(93)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(93) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initial_CP_1047_elements(93) is bound as output of CP function.
    -- CP-element group 94:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	89 
    -- CP-element group 94: 	108 
    -- CP-element group 94: 	112 
    -- CP-element group 94: 	132 
    -- CP-element group 94: marked-successors 
    -- CP-element group 94: 	90 
    -- CP-element group 94: 	92 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/aggregated_phi_update_ack
      -- CP-element group 94: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/phi_stmt_304_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/phi_stmt_304_update_completed__ps
      -- 
    -- logger for CP element group initial_CP_1047_elements(94)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(94)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(94) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initial_CP_1047_elements(94) is bound as output of CP function.
    -- CP-element group 95:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	86 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/phi_stmt_304_loopback_trigger
      -- 
    -- logger for CP element group initial_CP_1047_elements(95)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(95)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(95) fired."); 
        -- 
      end if; --
    end process; 
    initial_CP_1047_elements(95) <= initial_CP_1047_elements(86);
    -- CP-element group 96:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/phi_stmt_304_loopback_sample_req
      -- CP-element group 96: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/phi_stmt_304_loopback_sample_req_ps
      -- 
    -- logger for CP element group initial_CP_1047_elements(96)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(96)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(96) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:phi_stmt_304_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_304_loopback_sample_req_1518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_304_loopback_sample_req_1518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(96), ack => phi_stmt_304_req_1); -- 
    -- Element group initial_CP_1047_elements(96) is bound as output of CP function.
    -- CP-element group 97:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	87 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/phi_stmt_304_entry_trigger
      -- 
    -- logger for CP element group initial_CP_1047_elements(97)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(97)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(97) fired."); 
        -- 
      end if; --
    end process; 
    initial_CP_1047_elements(97) <= initial_CP_1047_elements(87);
    -- CP-element group 98:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/phi_stmt_304_entry_sample_req
      -- CP-element group 98: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/phi_stmt_304_entry_sample_req_ps
      -- 
    -- logger for CP element group initial_CP_1047_elements(98)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(98)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(98) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:phi_stmt_304_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_304_entry_sample_req_1521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_304_entry_sample_req_1521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(98), ack => phi_stmt_304_req_0); -- 
    -- Element group initial_CP_1047_elements(98) is bound as output of CP function.
    -- CP-element group 99:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/phi_stmt_304_phi_mux_ack
      -- CP-element group 99: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/phi_stmt_304_phi_mux_ack_ps
      -- 
    -- logger for CP element group initial_CP_1047_elements(99)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(99)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(99) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:phi_stmt_304_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_304_phi_mux_ack_1524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_304_ack_0, ack => initial_CP_1047_elements(99)); -- 
    -- CP-element group 100:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (4) 
      -- CP-element group 100: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_307_sample_start__ps
      -- CP-element group 100: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_307_sample_completed__ps
      -- CP-element group 100: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_307_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_307_sample_completed_
      -- 
    -- logger for CP element group initial_CP_1047_elements(100)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(100)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(100) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initial_CP_1047_elements(100) is bound as output of CP function.
    -- CP-element group 101:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_307_update_start__ps
      -- CP-element group 101: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_307_update_start_
      -- 
    -- logger for CP element group initial_CP_1047_elements(101)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(101)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(101) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initial_CP_1047_elements(101) is bound as output of CP function.
    -- CP-element group 102:  join  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	103 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_307_update_completed__ps
      -- 
    -- logger for CP element group initial_CP_1047_elements(102)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(102)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(102) fired."); 
        -- 
      end if; --
    end process; 
    initial_CP_1047_elements(102) <= initial_CP_1047_elements(103);
    -- CP-element group 103:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	102 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_307_update_completed_
      -- 
    -- logger for CP element group initial_CP_1047_elements(103)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(103)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(103) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initial_CP_1047_elements(103) is a control-delay.
    cp_element_103_delay: control_delay_element  generic map(name => " 103_delay", delay_value => 1)  port map(req => initial_CP_1047_elements(101), ack => initial_CP_1047_elements(103), clk => clk, reset =>reset);
    -- CP-element group 104:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (4) 
      -- CP-element group 104: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/R_NM_308_sample_start__ps
      -- CP-element group 104: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/R_NM_308_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/R_NM_308_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/R_NM_308_Sample/req
      -- 
    -- logger for CP element group initial_CP_1047_elements(104)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(104)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(104) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:NM_335_308_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(104), ack => NM_335_308_buf_req_0); -- 
    -- Element group initial_CP_1047_elements(104) is bound as output of CP function.
    -- CP-element group 105:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/R_NM_308_update_start__ps
      -- CP-element group 105: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/R_NM_308_update_start_
      -- CP-element group 105: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/R_NM_308_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/R_NM_308_Update/req
      -- 
    -- logger for CP element group initial_CP_1047_elements(105)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(105)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(105) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:NM_335_308_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(105), ack => NM_335_308_buf_req_1); -- 
    -- Element group initial_CP_1047_elements(105) is bound as output of CP function.
    -- CP-element group 106:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (4) 
      -- CP-element group 106: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/R_NM_308_sample_completed__ps
      -- CP-element group 106: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/R_NM_308_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/R_NM_308_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/R_NM_308_Sample/ack
      -- 
    -- logger for CP element group initial_CP_1047_elements(106)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(106)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(106) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:NM_335_308_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NM_335_308_buf_ack_0, ack => initial_CP_1047_elements(106)); -- 
    -- CP-element group 107:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (4) 
      -- CP-element group 107: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/R_NM_308_update_completed__ps
      -- CP-element group 107: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/R_NM_308_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/R_NM_308_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/R_NM_308_Update/ack
      -- 
    -- logger for CP element group initial_CP_1047_elements(107)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(107)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(107) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:NM_335_308_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NM_335_308_buf_ack_1, ack => initial_CP_1047_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	94 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	110 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_312_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_312_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_312_Sample/rr
      -- 
    -- logger for CP element group initial_CP_1047_elements(108)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(108)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(108) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:type_cast_312_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(108), ack => type_cast_312_inst_req_0); -- 
    initial_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "initial_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(94) & initial_CP_1047_elements(110);
      gj_initial_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	111 
    -- CP-element group 109: 	126 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_312_update_start_
      -- CP-element group 109: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_312_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_312_Update/cr
      -- 
    -- logger for CP element group initial_CP_1047_elements(109)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(109)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(109) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:type_cast_312_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(109), ack => type_cast_312_inst_req_1); -- 
    initial_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "initial_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(111) & initial_CP_1047_elements(126);
      gj_initial_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: marked-successors 
    -- CP-element group 110: 	92 
    -- CP-element group 110: 	108 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_312_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_312_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_312_Sample/ra
      -- 
    -- logger for CP element group initial_CP_1047_elements(110)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(110)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(110) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:type_cast_312_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_312_inst_ack_0, ack => initial_CP_1047_elements(110)); -- 
    -- CP-element group 111:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	124 
    -- CP-element group 111: marked-successors 
    -- CP-element group 111: 	109 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_312_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_312_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_312_Update/ca
      -- 
    -- logger for CP element group initial_CP_1047_elements(111)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(111)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(111) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:type_cast_312_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_312_inst_ack_1, ack => initial_CP_1047_elements(111)); -- 
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	94 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	114 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_316_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_316_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_316_Sample/req
      -- 
    -- logger for CP element group initial_CP_1047_elements(112)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(112)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(112) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:W_M_279_delayed_4_0_314_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(112), ack => W_M_279_delayed_4_0_314_inst_req_0); -- 
    initial_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "initial_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(94) & initial_CP_1047_elements(114);
      gj_initial_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	115 
    -- CP-element group 113: 	122 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_316_update_start_
      -- CP-element group 113: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_316_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_316_Update/req
      -- 
    -- logger for CP element group initial_CP_1047_elements(113)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(113)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(113) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:W_M_279_delayed_4_0_314_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(113), ack => W_M_279_delayed_4_0_314_inst_req_1); -- 
    initial_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "initial_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(115) & initial_CP_1047_elements(122);
      gj_initial_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: marked-successors 
    -- CP-element group 114: 	92 
    -- CP-element group 114: 	112 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_316_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_316_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_316_Sample/ack
      -- 
    -- logger for CP element group initial_CP_1047_elements(114)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(114)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(114) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:W_M_279_delayed_4_0_314_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_M_279_delayed_4_0_314_inst_ack_0, ack => initial_CP_1047_elements(114)); -- 
    -- CP-element group 115:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	113 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_316_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_316_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_316_Update/ack
      -- 
    -- logger for CP element group initial_CP_1047_elements(115)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(115)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(115) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:W_M_279_delayed_4_0_314_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_M_279_delayed_4_0_314_inst_ack_1, ack => initial_CP_1047_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: 	121 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	122 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	122 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_321_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_321_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_321_Sample/rr
      -- 
    -- logger for CP element group initial_CP_1047_elements(116)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(116)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(116) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:type_cast_321_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(116), ack => type_cast_321_inst_req_0); -- 
    initial_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "initial_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initial_CP_1047_elements(115) & initial_CP_1047_elements(121) & initial_CP_1047_elements(122);
      gj_initial_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	123 
    -- CP-element group 117: 	130 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	123 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_321_update_start_
      -- CP-element group 117: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_321_Update/$entry
      -- CP-element group 117: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_321_Update/cr
      -- 
    -- logger for CP element group initial_CP_1047_elements(117)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(117)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(117) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:type_cast_321_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(117), ack => type_cast_321_inst_req_1); -- 
    initial_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "initial_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(123) & initial_CP_1047_elements(130);
      gj_initial_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	88 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	120 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_Sample/word_access_start/$entry
      -- CP-element group 118: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_Sample/word_access_start/word_0/$entry
      -- CP-element group 118: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initial_CP_1047_elements(118)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(118)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(118) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:LOAD_ZJ_318_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(118), ack => LOAD_ZJ_318_load_0_req_0); -- 
    initial_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "initial_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(88) & initial_CP_1047_elements(120);
      gj_initial_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	121 
    -- CP-element group 119: 	122 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_update_start_
      -- CP-element group 119: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_Update/word_access_complete/$entry
      -- CP-element group 119: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_Update/word_access_complete/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group initial_CP_1047_elements(119)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(119)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(119) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:LOAD_ZJ_318_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(119), ack => LOAD_ZJ_318_load_0_req_1); -- 
    initial_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "initial_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(121) & initial_CP_1047_elements(122);
      gj_initial_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: marked-successors 
    -- CP-element group 120: 	118 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_sample_completed_
      -- CP-element group 120: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_Sample/word_access_start/$exit
      -- CP-element group 120: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_Sample/word_access_start/word_0/$exit
      -- CP-element group 120: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initial_CP_1047_elements(120)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(120)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(120) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:LOAD_ZJ_318_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ZJ_318_load_0_ack_0, ack => initial_CP_1047_elements(120)); -- 
    -- CP-element group 121:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	116 
    -- CP-element group 121: marked-successors 
    -- CP-element group 121: 	119 
    -- CP-element group 121:  members (9) 
      -- CP-element group 121: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_Update/word_access_complete/$exit
      -- CP-element group 121: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_Update/word_access_complete/word_0/$exit
      -- CP-element group 121: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_Update/word_access_complete/word_0/ca
      -- CP-element group 121: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_Update/LOAD_ZJ_318_Merge/$entry
      -- CP-element group 121: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_Update/LOAD_ZJ_318_Merge/$exit
      -- CP-element group 121: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_Update/LOAD_ZJ_318_Merge/merge_req
      -- CP-element group 121: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/LOAD_ZJ_318_Update/LOAD_ZJ_318_Merge/merge_ack
      -- 
    -- logger for CP element group initial_CP_1047_elements(121)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(121)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(121) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:LOAD_ZJ_318_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ZJ_318_load_0_ack_1, ack => initial_CP_1047_elements(121)); -- 
    -- CP-element group 122:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	116 
    -- CP-element group 122: successors 
    -- CP-element group 122: marked-successors 
    -- CP-element group 122: 	113 
    -- CP-element group 122: 	116 
    -- CP-element group 122: 	119 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_321_sample_completed_
      -- CP-element group 122: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_321_Sample/$exit
      -- CP-element group 122: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_321_Sample/ra
      -- 
    -- logger for CP element group initial_CP_1047_elements(122)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(122)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(122) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:type_cast_321_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_321_inst_ack_0, ack => initial_CP_1047_elements(122)); -- 
    -- CP-element group 123:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	117 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	128 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	117 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_321_update_completed_
      -- CP-element group 123: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_321_Update/$exit
      -- CP-element group 123: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/type_cast_321_Update/ca
      -- 
    -- logger for CP element group initial_CP_1047_elements(123)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(123)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(123) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:type_cast_321_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_321_inst_ack_1, ack => initial_CP_1047_elements(123)); -- 
    -- CP-element group 124:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	111 
    -- CP-element group 124: marked-predecessors 
    -- CP-element group 124: 	126 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_325_sample_start_
      -- CP-element group 124: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_325_Sample/$entry
      -- CP-element group 124: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_325_Sample/req
      -- 
    -- logger for CP element group initial_CP_1047_elements(124)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(124)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(124) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:W_wdata_285_delayed_4_0_323_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(124), ack => W_wdata_285_delayed_4_0_323_inst_req_0); -- 
    initial_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "initial_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(111) & initial_CP_1047_elements(126);
      gj_initial_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: marked-predecessors 
    -- CP-element group 125: 	127 
    -- CP-element group 125: 	130 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_325_update_start_
      -- CP-element group 125: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_325_Update/$entry
      -- CP-element group 125: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_325_Update/req
      -- 
    -- logger for CP element group initial_CP_1047_elements(125)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(125)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(125) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:W_wdata_285_delayed_4_0_323_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(125), ack => W_wdata_285_delayed_4_0_323_inst_req_1); -- 
    initial_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "initial_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(127) & initial_CP_1047_elements(130);
      gj_initial_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126: marked-successors 
    -- CP-element group 126: 	109 
    -- CP-element group 126: 	124 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_325_sample_completed_
      -- CP-element group 126: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_325_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_325_Sample/ack
      -- 
    -- logger for CP element group initial_CP_1047_elements(126)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(126)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(126) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:W_wdata_285_delayed_4_0_323_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_285_delayed_4_0_323_inst_ack_0, ack => initial_CP_1047_elements(126)); -- 
    -- CP-element group 127:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	125 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_325_update_completed_
      -- CP-element group 127: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_325_Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/assign_stmt_325_Update/ack
      -- 
    -- logger for CP element group initial_CP_1047_elements(127)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(127)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(127) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:W_wdata_285_delayed_4_0_323_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_285_delayed_4_0_323_inst_ack_1, ack => initial_CP_1047_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	123 
    -- CP-element group 128: 	127 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	130 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/call_stmt_330_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/call_stmt_330_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/call_stmt_330_Sample/crr
      -- 
    -- logger for CP element group initial_CP_1047_elements(128)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(128)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(128) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:call_stmt_330_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(128), ack => call_stmt_330_call_req_0); -- 
    initial_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "initial_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initial_CP_1047_elements(123) & initial_CP_1047_elements(127) & initial_CP_1047_elements(130);
      gj_initial_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	131 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/call_stmt_330_update_start_
      -- CP-element group 129: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/call_stmt_330_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/call_stmt_330_Update/ccr
      -- 
    -- logger for CP element group initial_CP_1047_elements(129)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(129)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(129) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:call_stmt_330_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_1654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(129), ack => call_stmt_330_call_req_1); -- 
    initial_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "initial_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= initial_CP_1047_elements(131);
      gj_initial_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: marked-successors 
    -- CP-element group 130: 	117 
    -- CP-element group 130: 	125 
    -- CP-element group 130: 	128 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/call_stmt_330_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/call_stmt_330_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/call_stmt_330_Sample/cra
      -- 
    -- logger for CP element group initial_CP_1047_elements(130)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(130)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(130) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:call_stmt_330_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_330_call_ack_0, ack => initial_CP_1047_elements(130)); -- 
    -- CP-element group 131:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	85 
    -- CP-element group 131: marked-successors 
    -- CP-element group 131: 	129 
    -- CP-element group 131:  members (4) 
      -- CP-element group 131: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/$exit
      -- CP-element group 131: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/call_stmt_330_update_completed_
      -- CP-element group 131: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/call_stmt_330_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/call_stmt_330_Update/cca
      -- 
    -- logger for CP element group initial_CP_1047_elements(131)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(131)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(131) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:call_stmt_330_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_330_call_ack_1, ack => initial_CP_1047_elements(131)); -- 
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	94 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/ADD_u12_u12_334_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/ADD_u12_u12_334_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/ADD_u12_u12_334_Sample/rr
      -- 
    -- logger for CP element group initial_CP_1047_elements(132)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(132)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(132) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:ADD_u12_u12_334_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(132), ack => ADD_u12_u12_334_inst_req_0); -- 
    initial_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "initial_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(94) & initial_CP_1047_elements(134);
      gj_initial_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	93 
    -- CP-element group 133: marked-predecessors 
    -- CP-element group 133: 	135 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	135 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/ADD_u12_u12_334_update_start_
      -- CP-element group 133: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/ADD_u12_u12_334_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/ADD_u12_u12_334_Update/cr
      -- 
    -- logger for CP element group initial_CP_1047_elements(133)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(133)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(133) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:ADD_u12_u12_334_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initial_CP_1047_elements(133), ack => ADD_u12_u12_334_inst_req_1); -- 
    initial_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "initial_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initial_CP_1047_elements(93) & initial_CP_1047_elements(135);
      gj_initial_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initial_CP_1047_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	92 
    -- CP-element group 134: 	132 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/ADD_u12_u12_334_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/ADD_u12_u12_334_Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/ADD_u12_u12_334_Sample/ra
      -- 
    -- logger for CP element group initial_CP_1047_elements(134)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(134)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(134) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:ADD_u12_u12_334_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_334_inst_ack_0, ack => initial_CP_1047_elements(134)); -- 
    -- CP-element group 135:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	89 
    -- CP-element group 135: marked-successors 
    -- CP-element group 135: 	91 
    -- CP-element group 135: 	133 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/ADD_u12_u12_334_update_completed_
      -- CP-element group 135: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/ADD_u12_u12_334_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/ADD_u12_u12_334_Update/ca
      -- 
    -- logger for CP element group initial_CP_1047_elements(135)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(135)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(135) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:ADD_u12_u12_334_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_334_inst_ack_1, ack => initial_CP_1047_elements(135)); -- 
    -- CP-element group 136:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	88 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	89 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_301/do_while_stmt_302/do_while_stmt_302_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group initial_CP_1047_elements(136)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(136)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(136) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initial_CP_1047_elements(136) is a control-delay.
    cp_element_136_delay: control_delay_element  generic map(name => " 136_delay", delay_value => 1)  port map(req => initial_CP_1047_elements(88), ack => initial_CP_1047_elements(136), clk => clk, reset =>reset);
    -- CP-element group 137:  transition  input  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	84 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (2) 
      -- CP-element group 137: 	 branch_block_stmt_301/do_while_stmt_302/loop_exit/ack
      -- CP-element group 137: 	 branch_block_stmt_301/do_while_stmt_302/loop_exit/$exit
      -- 
    -- logger for CP element group initial_CP_1047_elements(137)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(137)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(137) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:do_while_stmt_302_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_302_branch_ack_0, ack => initial_CP_1047_elements(137)); -- 
    -- CP-element group 138:  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	84 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (2) 
      -- CP-element group 138: 	 branch_block_stmt_301/do_while_stmt_302/loop_taken/ack
      -- CP-element group 138: 	 branch_block_stmt_301/do_while_stmt_302/loop_taken/$exit
      -- 
    -- logger for CP element group initial_CP_1047_elements(138)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(138)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(138) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:do_while_stmt_302_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_302_branch_ack_1, ack => initial_CP_1047_elements(138)); -- 
    -- CP-element group 139:  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	82 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	80 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_301/do_while_stmt_302/$exit
      -- 
    -- logger for CP element group initial_CP_1047_elements(139)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initial_CP_1047_elements(139)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initial:CP:initial_CP_1047_elements(139) fired."); 
        -- 
      end if; --
    end process; 
    initial_CP_1047_elements(139) <= initial_CP_1047_elements(82);
    initial_do_while_stmt_247_terminator_1348: loop_terminator -- 
      generic map (name => " initial_do_while_stmt_247_terminator_1348", max_iterations_in_flight =>7) 
      port map(loop_body_exit => initial_CP_1047_elements(13),loop_continue => initial_CP_1047_elements(66),loop_terminate => initial_CP_1047_elements(65),loop_back => initial_CP_1047_elements(11),loop_exit => initial_CP_1047_elements(10),clk => clk, reset => reset); -- 
    phi_stmt_249_phi_seq_1221_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= initial_CP_1047_elements(25);
      initial_CP_1047_elements(28)<= src_sample_reqs(0);
      src_sample_acks(0)  <= initial_CP_1047_elements(28);
      initial_CP_1047_elements(29)<= src_update_reqs(0);
      src_update_acks(0)  <= initial_CP_1047_elements(30);
      initial_CP_1047_elements(26) <= phi_mux_reqs(0);
      triggers(1)  <= initial_CP_1047_elements(23);
      initial_CP_1047_elements(32)<= src_sample_reqs(1);
      src_sample_acks(1)  <= initial_CP_1047_elements(34);
      initial_CP_1047_elements(33)<= src_update_reqs(1);
      src_update_acks(1)  <= initial_CP_1047_elements(35);
      initial_CP_1047_elements(24) <= phi_mux_reqs(1);
      phi_stmt_249_phi_seq_1221 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_249_phi_seq_1221") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => initial_CP_1047_elements(18), 
          phi_sample_ack => initial_CP_1047_elements(21), 
          phi_update_req => initial_CP_1047_elements(20), 
          phi_update_ack => initial_CP_1047_elements(22), 
          phi_mux_ack => initial_CP_1047_elements(27), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1173_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= initial_CP_1047_elements(14);
        preds(1)  <= initial_CP_1047_elements(15);
        entry_tmerge_1173 : transition_merge -- 
          generic map(name => " entry_tmerge_1173")
          port map (preds => preds, symbol_out => initial_CP_1047_elements(16));
          -- 
    end block;
    initial_do_while_stmt_302_terminator_1679: loop_terminator -- 
      generic map (name => " initial_do_while_stmt_302_terminator_1679", max_iterations_in_flight =>7) 
      port map(loop_body_exit => initial_CP_1047_elements(85),loop_continue => initial_CP_1047_elements(138),loop_terminate => initial_CP_1047_elements(137),loop_back => initial_CP_1047_elements(83),loop_exit => initial_CP_1047_elements(82),clk => clk, reset => reset); -- 
    phi_stmt_304_phi_seq_1552_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= initial_CP_1047_elements(97);
      initial_CP_1047_elements(100)<= src_sample_reqs(0);
      src_sample_acks(0)  <= initial_CP_1047_elements(100);
      initial_CP_1047_elements(101)<= src_update_reqs(0);
      src_update_acks(0)  <= initial_CP_1047_elements(102);
      initial_CP_1047_elements(98) <= phi_mux_reqs(0);
      triggers(1)  <= initial_CP_1047_elements(95);
      initial_CP_1047_elements(104)<= src_sample_reqs(1);
      src_sample_acks(1)  <= initial_CP_1047_elements(106);
      initial_CP_1047_elements(105)<= src_update_reqs(1);
      src_update_acks(1)  <= initial_CP_1047_elements(107);
      initial_CP_1047_elements(96) <= phi_mux_reqs(1);
      phi_stmt_304_phi_seq_1552 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_304_phi_seq_1552") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => initial_CP_1047_elements(90), 
          phi_sample_ack => initial_CP_1047_elements(93), 
          phi_update_req => initial_CP_1047_elements(92), 
          phi_update_ack => initial_CP_1047_elements(94), 
          phi_mux_ack => initial_CP_1047_elements(99), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1504_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= initial_CP_1047_elements(86);
        preds(1)  <= initial_CP_1047_elements(87);
        entry_tmerge_1504 : transition_merge -- 
          generic map(name => " entry_tmerge_1504")
          port map (preds => preds, symbol_out => initial_CP_1047_elements(88));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u12_u12_265_wire : std_logic_vector(11 downto 0);
    signal ADD_u12_u12_320_wire : std_logic_vector(11 downto 0);
    signal I_230_delayed_4_0_261 : std_logic_vector(11 downto 0);
    signal I_249 : std_logic_vector(11 downto 0);
    signal LOAD_ZJ_263_data_0 : std_logic_vector(11 downto 0);
    signal LOAD_ZJ_263_wire : std_logic_vector(11 downto 0);
    signal LOAD_ZJ_263_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_ZJ_318_data_0 : std_logic_vector(11 downto 0);
    signal LOAD_ZJ_318_wire : std_logic_vector(11 downto 0);
    signal LOAD_ZJ_318_word_address_0 : std_logic_vector(0 downto 0);
    signal MUL_u12_u12_244_wire : std_logic_vector(11 downto 0);
    signal M_279_delayed_4_0_316 : std_logic_vector(11 downto 0);
    signal M_304 : std_logic_vector(11 downto 0);
    signal NI_280 : std_logic_vector(11 downto 0);
    signal NI_280_253_buffered : std_logic_vector(11 downto 0);
    signal NM_335 : std_logic_vector(11 downto 0);
    signal NM_335_308_buffered : std_logic_vector(11 downto 0);
    signal STORE_ZJ_230_data_0 : std_logic_vector(11 downto 0);
    signal STORE_ZJ_230_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_ZJ_241_data_0 : std_logic_vector(11 downto 0);
    signal STORE_ZJ_241_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_ZJ_298_data_0 : std_logic_vector(11 downto 0);
    signal STORE_ZJ_298_word_address_0 : std_logic_vector(0 downto 0);
    signal ULT_u12_u1_284_wire : std_logic_vector(0 downto 0);
    signal ULT_u12_u1_294_wire : std_logic_vector(0 downto 0);
    signal ULT_u12_u1_339_wire : std_logic_vector(0 downto 0);
    signal YI_290 : std_logic_vector(11 downto 0);
    signal YI_290_239_buffered : std_logic_vector(11 downto 0);
    signal Y_235 : std_logic_vector(11 downto 0);
    signal addr_267 : std_logic_vector(11 downto 0);
    signal addr_322 : std_logic_vector(11 downto 0);
    signal konst_231_wire_constant : std_logic_vector(11 downto 0);
    signal konst_243_wire_constant : std_logic_vector(11 downto 0);
    signal konst_271_wire_constant : std_logic_vector(0 downto 0);
    signal konst_278_wire_constant : std_logic_vector(11 downto 0);
    signal konst_283_wire_constant : std_logic_vector(11 downto 0);
    signal konst_288_wire_constant : std_logic_vector(11 downto 0);
    signal konst_293_wire_constant : std_logic_vector(11 downto 0);
    signal konst_299_wire_constant : std_logic_vector(11 downto 0);
    signal konst_326_wire_constant : std_logic_vector(0 downto 0);
    signal konst_333_wire_constant : std_logic_vector(11 downto 0);
    signal konst_338_wire_constant : std_logic_vector(11 downto 0);
    signal rdata_275 : std_logic_vector(63 downto 0);
    signal rdata_330 : std_logic_vector(63 downto 0);
    signal type_cast_238_wire_constant : std_logic_vector(11 downto 0);
    signal type_cast_252_wire_constant : std_logic_vector(11 downto 0);
    signal type_cast_307_wire_constant : std_logic_vector(11 downto 0);
    signal wdata_236_delayed_4_0_270 : std_logic_vector(15 downto 0);
    signal wdata_258 : std_logic_vector(15 downto 0);
    signal wdata_285_delayed_4_0_325 : std_logic_vector(15 downto 0);
    signal wdata_313 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    LOAD_ZJ_263_word_address_0 <= "0";
    LOAD_ZJ_318_word_address_0 <= "0";
    STORE_ZJ_230_word_address_0 <= "0";
    STORE_ZJ_241_word_address_0 <= "0";
    STORE_ZJ_298_word_address_0 <= "0";
    konst_231_wire_constant <= "000000000000";
    konst_243_wire_constant <= "000010000000";
    konst_271_wire_constant <= "0";
    konst_278_wire_constant <= "000000000001";
    konst_283_wire_constant <= "000010000000";
    konst_288_wire_constant <= "000000000001";
    konst_293_wire_constant <= "000000001000";
    konst_299_wire_constant <= "010000000000";
    konst_326_wire_constant <= "0";
    konst_333_wire_constant <= "000000000001";
    konst_338_wire_constant <= "000000010000";
    type_cast_238_wire_constant <= "000000000000";
    type_cast_252_wire_constant <= "000000000000";
    type_cast_307_wire_constant <= "000000000000";
    -- logger for phi phi_stmt_235
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_235_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:initial:DP:phi_stmt_235:input-0 type_cast_238_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_238_wire_constant));
          --
        end if;
        if phi_stmt_235_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:initial:DP:phi_stmt_235:input-1 YI_290_239_buffered= " & Convert_SLV_To_Hex_String(YI_290_239_buffered));
          --
        end if;
        if phi_stmt_235_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:initial:DP:phi_stmt_235:sample-completed");
          --
        end if;
        if phi_stmt_235_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:initial:DP:phi_stmt_235:output Y_235= " & Convert_SLV_To_Hex_String(Y_235));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_235: Block -- phi operator 
      signal idata: std_logic_vector(23 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_238_wire_constant & YI_290_239_buffered;
      req <= phi_stmt_235_req_0 & phi_stmt_235_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_235",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 12) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_235_ack_0,
          idata => idata,
          odata => Y_235,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_235
    -- logger for phi phi_stmt_249
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_249_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:initial:DP:phi_stmt_249:input-0 type_cast_252_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_252_wire_constant));
          --
        end if;
        if phi_stmt_249_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:initial:DP:phi_stmt_249:input-1 NI_280_253_buffered= " & Convert_SLV_To_Hex_String(NI_280_253_buffered));
          --
        end if;
        if phi_stmt_249_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:initial:DP:phi_stmt_249:sample-completed");
          --
        end if;
        if phi_stmt_249_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:initial:DP:phi_stmt_249:output I_249= " & Convert_SLV_To_Hex_String(I_249));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_249: Block -- phi operator 
      signal idata: std_logic_vector(23 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_252_wire_constant & NI_280_253_buffered;
      req <= phi_stmt_249_req_0 & phi_stmt_249_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_249",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 12) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_249_ack_0,
          idata => idata,
          odata => I_249,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_249
    -- logger for phi phi_stmt_304
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_304_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:initial:DP:phi_stmt_304:input-0 type_cast_307_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_307_wire_constant));
          --
        end if;
        if phi_stmt_304_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:initial:DP:phi_stmt_304:input-1 NM_335_308_buffered= " & Convert_SLV_To_Hex_String(NM_335_308_buffered));
          --
        end if;
        if phi_stmt_304_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:initial:DP:phi_stmt_304:sample-completed");
          --
        end if;
        if phi_stmt_304_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:initial:DP:phi_stmt_304:output M_304= " & Convert_SLV_To_Hex_String(M_304));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_304: Block -- phi operator 
      signal idata: std_logic_vector(23 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_307_wire_constant & NM_335_308_buffered;
      req <= phi_stmt_304_req_0 & phi_stmt_304_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_304",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 12) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_304_ack_0,
          idata => idata,
          odata => M_304,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_304
    -- logger for split-operator NI_280_253_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if NI_280_253_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:NI_280_253_buf:started:   inputs: " & " NI_280 = "& Convert_SLV_To_Hex_String(NI_280));
          --
        end if; 
        if NI_280_253_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:NI_280_253_buf:finished:  outputs: " & " NI_280_253_buffered= "  & Convert_SLV_To_Hex_String(NI_280_253_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    NI_280_253_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= NI_280_253_buf_req_0;
      NI_280_253_buf_ack_0<= wack(0);
      rreq(0) <= NI_280_253_buf_req_1;
      NI_280_253_buf_ack_1<= rack(0);
      NI_280_253_buf : InterlockBuffer generic map ( -- 
        name => "NI_280_253_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => NI_280,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NI_280_253_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator NM_335_308_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if NM_335_308_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:NM_335_308_buf:started:   inputs: " & " NM_335 = "& Convert_SLV_To_Hex_String(NM_335));
          --
        end if; 
        if NM_335_308_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:NM_335_308_buf:finished:  outputs: " & " NM_335_308_buffered= "  & Convert_SLV_To_Hex_String(NM_335_308_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    NM_335_308_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= NM_335_308_buf_req_0;
      NM_335_308_buf_ack_0<= wack(0);
      rreq(0) <= NM_335_308_buf_req_1;
      NM_335_308_buf_ack_1<= rack(0);
      NM_335_308_buf : InterlockBuffer generic map ( -- 
        name => "NM_335_308_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => NM_335,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NM_335_308_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_I_230_delayed_4_0_259_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_I_230_delayed_4_0_259_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:W_I_230_delayed_4_0_259_inst:started:   inputs: " & " I_249 = "& Convert_SLV_To_Hex_String(I_249));
          --
        end if; 
        if W_I_230_delayed_4_0_259_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:W_I_230_delayed_4_0_259_inst:finished:  outputs: " & " I_230_delayed_4_0_261= "  & Convert_SLV_To_Hex_String(I_230_delayed_4_0_261));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_I_230_delayed_4_0_259_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_I_230_delayed_4_0_259_inst_req_0;
      W_I_230_delayed_4_0_259_inst_ack_0<= wack(0);
      rreq(0) <= W_I_230_delayed_4_0_259_inst_req_1;
      W_I_230_delayed_4_0_259_inst_ack_1<= rack(0);
      W_I_230_delayed_4_0_259_inst : InterlockBuffer generic map ( -- 
        name => "W_I_230_delayed_4_0_259_inst",
        buffer_size => 4,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => I_249,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => I_230_delayed_4_0_261,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_M_279_delayed_4_0_314_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_M_279_delayed_4_0_314_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:W_M_279_delayed_4_0_314_inst:started:   inputs: " & " M_304 = "& Convert_SLV_To_Hex_String(M_304));
          --
        end if; 
        if W_M_279_delayed_4_0_314_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:W_M_279_delayed_4_0_314_inst:finished:  outputs: " & " M_279_delayed_4_0_316= "  & Convert_SLV_To_Hex_String(M_279_delayed_4_0_316));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_M_279_delayed_4_0_314_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_M_279_delayed_4_0_314_inst_req_0;
      W_M_279_delayed_4_0_314_inst_ack_0<= wack(0);
      rreq(0) <= W_M_279_delayed_4_0_314_inst_req_1;
      W_M_279_delayed_4_0_314_inst_ack_1<= rack(0);
      W_M_279_delayed_4_0_314_inst : InterlockBuffer generic map ( -- 
        name => "W_M_279_delayed_4_0_314_inst",
        buffer_size => 4,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => M_304,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => M_279_delayed_4_0_316,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_wdata_236_delayed_4_0_268_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_wdata_236_delayed_4_0_268_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:W_wdata_236_delayed_4_0_268_inst:started:   inputs: " & " wdata_258 = "& Convert_SLV_To_Hex_String(wdata_258));
          --
        end if; 
        if W_wdata_236_delayed_4_0_268_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:W_wdata_236_delayed_4_0_268_inst:finished:  outputs: " & " wdata_236_delayed_4_0_270= "  & Convert_SLV_To_Hex_String(wdata_236_delayed_4_0_270));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_wdata_236_delayed_4_0_268_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_wdata_236_delayed_4_0_268_inst_req_0;
      W_wdata_236_delayed_4_0_268_inst_ack_0<= wack(0);
      rreq(0) <= W_wdata_236_delayed_4_0_268_inst_req_1;
      W_wdata_236_delayed_4_0_268_inst_ack_1<= rack(0);
      W_wdata_236_delayed_4_0_268_inst : InterlockBuffer generic map ( -- 
        name => "W_wdata_236_delayed_4_0_268_inst",
        buffer_size => 4,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => wdata_258,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => wdata_236_delayed_4_0_270,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_wdata_285_delayed_4_0_323_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_wdata_285_delayed_4_0_323_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:W_wdata_285_delayed_4_0_323_inst:started:   inputs: " & " wdata_313 = "& Convert_SLV_To_Hex_String(wdata_313));
          --
        end if; 
        if W_wdata_285_delayed_4_0_323_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:W_wdata_285_delayed_4_0_323_inst:finished:  outputs: " & " wdata_285_delayed_4_0_325= "  & Convert_SLV_To_Hex_String(wdata_285_delayed_4_0_325));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_wdata_285_delayed_4_0_323_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_wdata_285_delayed_4_0_323_inst_req_0;
      W_wdata_285_delayed_4_0_323_inst_ack_0<= wack(0);
      rreq(0) <= W_wdata_285_delayed_4_0_323_inst_req_1;
      W_wdata_285_delayed_4_0_323_inst_ack_1<= rack(0);
      W_wdata_285_delayed_4_0_323_inst : InterlockBuffer generic map ( -- 
        name => "W_wdata_285_delayed_4_0_323_inst",
        buffer_size => 4,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => wdata_313,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => wdata_285_delayed_4_0_325,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator YI_290_239_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if YI_290_239_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:YI_290_239_buf:started:   inputs: " & " YI_290 = "& Convert_SLV_To_Hex_String(YI_290));
          --
        end if; 
        if YI_290_239_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:YI_290_239_buf:finished:  outputs: " & " YI_290_239_buffered= "  & Convert_SLV_To_Hex_String(YI_290_239_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    YI_290_239_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= YI_290_239_buf_req_0;
      YI_290_239_buf_ack_0<= wack(0);
      rreq(0) <= YI_290_239_buf_req_1;
      YI_290_239_buf_ack_1<= rack(0);
      YI_290_239_buf : InterlockBuffer generic map ( -- 
        name => "YI_290_239_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => YI_290,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => YI_290_239_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_257_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_257_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:type_cast_257_inst:started:   inputs: " & " I_249 = "& Convert_SLV_To_Hex_String(I_249));
          --
        end if; 
        if type_cast_257_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:type_cast_257_inst:finished:  outputs: " & " wdata_258= "  & Convert_SLV_To_Hex_String(wdata_258));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_257_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_257_inst_req_0;
      type_cast_257_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_257_inst_req_1;
      type_cast_257_inst_ack_1<= rack(0);
      type_cast_257_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_257_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 12,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => I_249,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => wdata_258,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_266_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_266_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:type_cast_266_inst:started:   inputs: " & " ADD_u12_u12_265_wire = "& Convert_SLV_To_Hex_String(ADD_u12_u12_265_wire));
          --
        end if; 
        if type_cast_266_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:type_cast_266_inst:finished:  outputs: " & " addr_267= "  & Convert_SLV_To_Hex_String(addr_267));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_266_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_266_inst_req_0;
      type_cast_266_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_266_inst_req_1;
      type_cast_266_inst_ack_1<= rack(0);
      type_cast_266_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_266_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u12_u12_265_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => addr_267,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_312_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_312_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:type_cast_312_inst:started:   inputs: " & " M_304 = "& Convert_SLV_To_Hex_String(M_304));
          --
        end if; 
        if type_cast_312_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:type_cast_312_inst:finished:  outputs: " & " wdata_313= "  & Convert_SLV_To_Hex_String(wdata_313));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_312_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_312_inst_req_0;
      type_cast_312_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_312_inst_req_1;
      type_cast_312_inst_ack_1<= rack(0);
      type_cast_312_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_312_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 12,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => M_304,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => wdata_313,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_321_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_321_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:type_cast_321_inst:started:   inputs: " & " ADD_u12_u12_320_wire = "& Convert_SLV_To_Hex_String(ADD_u12_u12_320_wire));
          --
        end if; 
        if type_cast_321_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:type_cast_321_inst:finished:  outputs: " & " addr_322= "  & Convert_SLV_To_Hex_String(addr_322));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_321_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_321_inst_req_0;
      type_cast_321_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_321_inst_req_1;
      type_cast_321_inst_ack_1<= rack(0);
      type_cast_321_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_321_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u12_u12_320_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => addr_322,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for operator LOAD_ZJ_263_gather_scatter flow-through 
    process(LOAD_ZJ_263_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:LOAD_ZJ_263_gather_scatter:flowthrough  inputs: " & " LOAD_ZJ_263_data_0 = "& Convert_SLV_To_Hex_String(LOAD_ZJ_263_data_0) & "outputs: " & " LOAD_ZJ_263_wire= "  & Convert_SLV_To_Hex_String(LOAD_ZJ_263_wire));
      --
    end process; 
    -- equivalence LOAD_ZJ_263_gather_scatter
    process(LOAD_ZJ_263_data_0) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(11 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_ZJ_263_data_0;
      ov(11 downto 0) := iv;
      LOAD_ZJ_263_wire <= ov(11 downto 0);
      --
    end process;
    -- logger for operator LOAD_ZJ_318_gather_scatter flow-through 
    process(LOAD_ZJ_318_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:LOAD_ZJ_318_gather_scatter:flowthrough  inputs: " & " LOAD_ZJ_318_data_0 = "& Convert_SLV_To_Hex_String(LOAD_ZJ_318_data_0) & "outputs: " & " LOAD_ZJ_318_wire= "  & Convert_SLV_To_Hex_String(LOAD_ZJ_318_wire));
      --
    end process; 
    -- equivalence LOAD_ZJ_318_gather_scatter
    process(LOAD_ZJ_318_data_0) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(11 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_ZJ_318_data_0;
      ov(11 downto 0) := iv;
      LOAD_ZJ_318_wire <= ov(11 downto 0);
      --
    end process;
    -- logger for operator STORE_ZJ_230_gather_scatter flow-through 
    process(STORE_ZJ_230_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:STORE_ZJ_230_gather_scatter:flowthrough  inputs: " & " konst_231_wire_constant = "& Convert_SLV_To_Hex_String(konst_231_wire_constant) & "outputs: " & " STORE_ZJ_230_data_0= "  & Convert_SLV_To_Hex_String(STORE_ZJ_230_data_0));
      --
    end process; 
    -- equivalence STORE_ZJ_230_gather_scatter
    process(konst_231_wire_constant) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(11 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := konst_231_wire_constant;
      ov(11 downto 0) := iv;
      STORE_ZJ_230_data_0 <= ov(11 downto 0);
      --
    end process;
    -- logger for operator STORE_ZJ_241_gather_scatter flow-through 
    process(STORE_ZJ_241_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:STORE_ZJ_241_gather_scatter:flowthrough  inputs: " & " MUL_u12_u12_244_wire = "& Convert_SLV_To_Hex_String(MUL_u12_u12_244_wire) & "outputs: " & " STORE_ZJ_241_data_0= "  & Convert_SLV_To_Hex_String(STORE_ZJ_241_data_0));
      --
    end process; 
    -- equivalence STORE_ZJ_241_gather_scatter
    process(MUL_u12_u12_244_wire) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(11 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := MUL_u12_u12_244_wire;
      ov(11 downto 0) := iv;
      STORE_ZJ_241_data_0 <= ov(11 downto 0);
      --
    end process;
    -- logger for operator STORE_ZJ_298_gather_scatter flow-through 
    process(STORE_ZJ_298_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:STORE_ZJ_298_gather_scatter:flowthrough  inputs: " & " konst_299_wire_constant = "& Convert_SLV_To_Hex_String(konst_299_wire_constant) & "outputs: " & " STORE_ZJ_298_data_0= "  & Convert_SLV_To_Hex_String(STORE_ZJ_298_data_0));
      --
    end process; 
    -- equivalence STORE_ZJ_298_gather_scatter
    process(konst_299_wire_constant) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(11 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := konst_299_wire_constant;
      ov(11 downto 0) := iv;
      STORE_ZJ_298_data_0 <= ov(11 downto 0);
      --
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_247_branch_req_0," req0 do_while_stmt_247_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_247_branch_ack_0," ack0 do_while_stmt_247_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_247_branch_ack_1," ack1 do_while_stmt_247_branch");
    do_while_stmt_247_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u12_u1_284_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_247_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_247_branch_req_0,
          ack0 => do_while_stmt_247_branch_ack_0,
          ack1 => do_while_stmt_247_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_302_branch_req_0," req0 do_while_stmt_302_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_302_branch_ack_0," ack0 do_while_stmt_302_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_302_branch_ack_1," ack1 do_while_stmt_302_branch");
    do_while_stmt_302_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u12_u1_339_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_302_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_302_branch_req_0,
          ack0 => do_while_stmt_302_branch_ack_0,
          ack1 => do_while_stmt_302_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_291_branch_req_0," req0 if_stmt_291_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_291_branch_ack_0," ack0 if_stmt_291_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_291_branch_ack_1," ack1 if_stmt_291_branch");
    if_stmt_291_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u12_u1_294_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_291_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_291_branch_req_0,
          ack0 => if_stmt_291_branch_ack_0,
          ack1 => if_stmt_291_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator ADD_u12_u12_265_inst flow-through 
    process(ADD_u12_u12_265_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:ADD_u12_u12_265_inst:flowthrough inputs: " & " LOAD_ZJ_263_wire = "& Convert_SLV_To_Hex_String(LOAD_ZJ_263_wire) & " I_230_delayed_4_0_261 = "& Convert_SLV_To_Hex_String(I_230_delayed_4_0_261) & " outputs:" & " ADD_u12_u12_265_wire= "  & Convert_SLV_To_Hex_String(ADD_u12_u12_265_wire));
      --
    end process; 
    -- binary operator ADD_u12_u12_265_inst
    process(LOAD_ZJ_263_wire, I_230_delayed_4_0_261) -- 
      variable tmp_var : std_logic_vector(11 downto 0); -- 
    begin -- 
      ApIntAdd_proc(LOAD_ZJ_263_wire, I_230_delayed_4_0_261, tmp_var);
      ADD_u12_u12_265_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u12_u12_279_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_279_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:ADD_u12_u12_279_inst:started:   inputs: " & " I_249 = "& Convert_SLV_To_Hex_String(I_249) & " konst_278_wire_constant = "& Convert_SLV_To_Hex_String(konst_278_wire_constant));
          --
        end if; 
        if ADD_u12_u12_279_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:ADD_u12_u12_279_inst:finished:  outputs: " & " NI_280= "  & Convert_SLV_To_Hex_String(NI_280));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (1) : ADD_u12_u12_279_inst 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= I_249;
      NI_280 <= data_out(11 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u12_u12_279_inst_req_0;
      ADD_u12_u12_279_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_279_inst_req_1;
      ADD_u12_u12_279_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000000000001",
          constant_width => 12,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- logger for split-operator ADD_u12_u12_289_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_289_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:ADD_u12_u12_289_inst:started:   inputs: " & " Y_235 = "& Convert_SLV_To_Hex_String(Y_235) & " konst_288_wire_constant = "& Convert_SLV_To_Hex_String(konst_288_wire_constant));
          --
        end if; 
        if ADD_u12_u12_289_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:ADD_u12_u12_289_inst:finished:  outputs: " & " YI_290= "  & Convert_SLV_To_Hex_String(YI_290));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (2) : ADD_u12_u12_289_inst 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= Y_235;
      YI_290 <= data_out(11 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u12_u12_289_inst_req_0;
      ADD_u12_u12_289_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_289_inst_req_1;
      ADD_u12_u12_289_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_2_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000000000001",
          constant_width => 12,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- logger for split-operator ADD_u12_u12_320_inst flow-through 
    process(ADD_u12_u12_320_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:ADD_u12_u12_320_inst:flowthrough inputs: " & " LOAD_ZJ_318_wire = "& Convert_SLV_To_Hex_String(LOAD_ZJ_318_wire) & " M_279_delayed_4_0_316 = "& Convert_SLV_To_Hex_String(M_279_delayed_4_0_316) & " outputs:" & " ADD_u12_u12_320_wire= "  & Convert_SLV_To_Hex_String(ADD_u12_u12_320_wire));
      --
    end process; 
    -- binary operator ADD_u12_u12_320_inst
    process(LOAD_ZJ_318_wire, M_279_delayed_4_0_316) -- 
      variable tmp_var : std_logic_vector(11 downto 0); -- 
    begin -- 
      ApIntAdd_proc(LOAD_ZJ_318_wire, M_279_delayed_4_0_316, tmp_var);
      ADD_u12_u12_320_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u12_u12_334_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_334_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:ADD_u12_u12_334_inst:started:   inputs: " & " M_304 = "& Convert_SLV_To_Hex_String(M_304) & " konst_333_wire_constant = "& Convert_SLV_To_Hex_String(konst_333_wire_constant));
          --
        end if; 
        if ADD_u12_u12_334_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:ADD_u12_u12_334_inst:finished:  outputs: " & " NM_335= "  & Convert_SLV_To_Hex_String(NM_335));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (4) : ADD_u12_u12_334_inst 
    ApIntAdd_group_4: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= M_304;
      NM_335 <= data_out(11 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u12_u12_334_inst_req_0;
      ADD_u12_u12_334_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_334_inst_req_1;
      ADD_u12_u12_334_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_4_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000000000001",
          constant_width => 12,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- logger for split-operator MUL_u12_u12_244_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if MUL_u12_u12_244_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:MUL_u12_u12_244_inst:started:   inputs: " & " Y_235 = "& Convert_SLV_To_Hex_String(Y_235) & " konst_243_wire_constant = "& Convert_SLV_To_Hex_String(konst_243_wire_constant));
          --
        end if; 
        if MUL_u12_u12_244_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:MUL_u12_u12_244_inst:finished:  outputs: " & " MUL_u12_u12_244_wire= "  & Convert_SLV_To_Hex_String(MUL_u12_u12_244_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (5) : MUL_u12_u12_244_inst 
    ApIntMul_group_5: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= Y_235;
      MUL_u12_u12_244_wire <= data_out(11 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= MUL_u12_u12_244_inst_req_0;
      MUL_u12_u12_244_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= MUL_u12_u12_244_inst_req_1;
      MUL_u12_u12_244_inst_ack_1 <= ackR_unguarded(0);
      ApIntMul_group_5_gI: SplitGuardInterface generic map(name => "ApIntMul_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          name => "ApIntMul_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000010000000",
          constant_width => 12,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- logger for split-operator ULT_u12_u1_284_inst flow-through 
    process(ULT_u12_u1_284_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:ULT_u12_u1_284_inst:flowthrough inputs: " & " NI_280 = "& Convert_SLV_To_Hex_String(NI_280) & " konst_283_wire_constant = "& Convert_SLV_To_Hex_String(konst_283_wire_constant) & " outputs:" & " ULT_u12_u1_284_wire= "  & Convert_SLV_To_Hex_String(ULT_u12_u1_284_wire));
      --
    end process; 
    -- binary operator ULT_u12_u1_284_inst
    process(NI_280) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(NI_280, konst_283_wire_constant, tmp_var);
      ULT_u12_u1_284_wire <= tmp_var; --
    end process;
    -- logger for split-operator ULT_u12_u1_294_inst flow-through 
    process(ULT_u12_u1_294_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:ULT_u12_u1_294_inst:flowthrough inputs: " & " YI_290 = "& Convert_SLV_To_Hex_String(YI_290) & " konst_293_wire_constant = "& Convert_SLV_To_Hex_String(konst_293_wire_constant) & " outputs:" & " ULT_u12_u1_294_wire= "  & Convert_SLV_To_Hex_String(ULT_u12_u1_294_wire));
      --
    end process; 
    -- binary operator ULT_u12_u1_294_inst
    process(YI_290) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(YI_290, konst_293_wire_constant, tmp_var);
      ULT_u12_u1_294_wire <= tmp_var; --
    end process;
    -- logger for split-operator ULT_u12_u1_339_inst flow-through 
    process(ULT_u12_u1_339_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:ULT_u12_u1_339_inst:flowthrough inputs: " & " NM_335 = "& Convert_SLV_To_Hex_String(NM_335) & " konst_338_wire_constant = "& Convert_SLV_To_Hex_String(konst_338_wire_constant) & " outputs:" & " ULT_u12_u1_339_wire= "  & Convert_SLV_To_Hex_String(ULT_u12_u1_339_wire));
      --
    end process; 
    -- binary operator ULT_u12_u1_339_inst
    process(NM_335) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(NM_335, konst_338_wire_constant, tmp_var);
      ULT_u12_u1_339_wire <= tmp_var; --
    end process;
    -- logger for split-operator LOAD_ZJ_263_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if LOAD_ZJ_263_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:LOAD_ZJ_263_load_0:started:   inputs: " & " LOAD_ZJ_263_word_address_0 = "& Convert_SLV_To_Hex_String(LOAD_ZJ_263_word_address_0));
          --
        end if; 
        if LOAD_ZJ_263_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:LOAD_ZJ_263_load_0:finished:  outputs: " & " LOAD_ZJ_263_data_0= "  & Convert_SLV_To_Hex_String(LOAD_ZJ_263_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator LOAD_ZJ_318_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if LOAD_ZJ_318_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:LOAD_ZJ_318_load_0:started:   inputs: " & " LOAD_ZJ_318_word_address_0 = "& Convert_SLV_To_Hex_String(LOAD_ZJ_318_word_address_0));
          --
        end if; 
        if LOAD_ZJ_318_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:LOAD_ZJ_318_load_0:finished:  outputs: " & " LOAD_ZJ_318_data_0= "  & Convert_SLV_To_Hex_String(LOAD_ZJ_318_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (0) : LOAD_ZJ_263_load_0 LOAD_ZJ_318_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 5, 1 => 5);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        LOAD_ZJ_263_load_0_req_0,
        LOAD_ZJ_263_load_0_ack_0,
        LOAD_ZJ_263_load_0_req_1,
        LOAD_ZJ_263_load_0_ack_1,
        "LOAD_ZJ_263_load_0",
        "memory_space_1" ,
        LOAD_ZJ_263_data_0,
        LOAD_ZJ_263_word_address_0,
        "LOAD_ZJ_263_data_0",
        "LOAD_ZJ_263_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        LOAD_ZJ_318_load_0_req_0,
        LOAD_ZJ_318_load_0_ack_0,
        LOAD_ZJ_318_load_0_req_1,
        LOAD_ZJ_318_load_0_ack_1,
        "LOAD_ZJ_318_load_0",
        "memory_space_1" ,
        LOAD_ZJ_318_data_0,
        LOAD_ZJ_318_word_address_0,
        "LOAD_ZJ_318_data_0",
        "LOAD_ZJ_318_word_address_0" -- 
      );
      reqL_unguarded(1) <= LOAD_ZJ_263_load_0_req_0;
      reqL_unguarded(0) <= LOAD_ZJ_318_load_0_req_0;
      LOAD_ZJ_263_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_ZJ_318_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= LOAD_ZJ_263_load_0_req_1;
      reqR_unguarded(0) <= LOAD_ZJ_318_load_0_req_1;
      LOAD_ZJ_263_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_ZJ_318_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_ZJ_263_word_address_0 & LOAD_ZJ_318_word_address_0;
      LOAD_ZJ_263_data_0 <= data_out(23 downto 12);
      LOAD_ZJ_318_data_0 <= data_out(11 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(0 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 12,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(11 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logger for split-operator STORE_ZJ_298_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if STORE_ZJ_298_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:STORE_ZJ_298_store_0:started:   inputs: " & " STORE_ZJ_298_word_address_0 = "& Convert_SLV_To_Hex_String(STORE_ZJ_298_word_address_0) & " STORE_ZJ_298_data_0 = "& Convert_SLV_To_Hex_String(STORE_ZJ_298_data_0));
          --
        end if; 
        if STORE_ZJ_298_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:STORE_ZJ_298_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator STORE_ZJ_230_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if STORE_ZJ_230_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:STORE_ZJ_230_store_0:started:   inputs: " & " STORE_ZJ_230_word_address_0 = "& Convert_SLV_To_Hex_String(STORE_ZJ_230_word_address_0) & " STORE_ZJ_230_data_0 = "& Convert_SLV_To_Hex_String(STORE_ZJ_230_data_0));
          --
        end if; 
        if STORE_ZJ_230_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:STORE_ZJ_230_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator STORE_ZJ_241_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if STORE_ZJ_241_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:STORE_ZJ_241_store_0:started:   inputs: " & " STORE_ZJ_241_word_address_0 = "& Convert_SLV_To_Hex_String(STORE_ZJ_241_word_address_0) & " STORE_ZJ_241_data_0 = "& Convert_SLV_To_Hex_String(STORE_ZJ_241_data_0));
          --
        end if; 
        if STORE_ZJ_241_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:STORE_ZJ_241_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      STORE_ZJ_298_store_0_req_0,
      STORE_ZJ_298_store_0_ack_0,
      STORE_ZJ_298_store_0_req_1,
      STORE_ZJ_298_store_0_ack_1,
      "STORE_ZJ_298_store_0",
      "memory_space_1" ,
      STORE_ZJ_298_data_0,
      STORE_ZJ_298_word_address_0,
      "STORE_ZJ_298_data_0",
      "STORE_ZJ_298_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      STORE_ZJ_230_store_0_req_0,
      STORE_ZJ_230_store_0_ack_0,
      STORE_ZJ_230_store_0_req_1,
      STORE_ZJ_230_store_0_ack_1,
      "STORE_ZJ_230_store_0",
      "memory_space_1" ,
      STORE_ZJ_230_data_0,
      STORE_ZJ_230_word_address_0,
      "STORE_ZJ_230_data_0",
      "STORE_ZJ_230_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      STORE_ZJ_241_store_0_req_0,
      STORE_ZJ_241_store_0_ack_0,
      STORE_ZJ_241_store_0_req_1,
      STORE_ZJ_241_store_0_ack_1,
      "STORE_ZJ_241_store_0",
      "memory_space_1" ,
      STORE_ZJ_241_data_0,
      STORE_ZJ_241_word_address_0,
      "STORE_ZJ_241_data_0",
      "STORE_ZJ_241_word_address_0" -- 
    );
    -- shared store operator group (0) : STORE_ZJ_298_store_0 STORE_ZJ_230_store_0 STORE_ZJ_241_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(2 downto 0);
      signal data_in: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= STORE_ZJ_298_store_0_req_0;
      reqL_unguarded(1) <= STORE_ZJ_230_store_0_req_0;
      reqL_unguarded(0) <= STORE_ZJ_241_store_0_req_0;
      STORE_ZJ_298_store_0_ack_0 <= ackL_unguarded(2);
      STORE_ZJ_230_store_0_ack_0 <= ackL_unguarded(1);
      STORE_ZJ_241_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= STORE_ZJ_298_store_0_req_1;
      reqR_unguarded(1) <= STORE_ZJ_230_store_0_req_1;
      reqR_unguarded(0) <= STORE_ZJ_241_store_0_req_1;
      STORE_ZJ_298_store_0_ack_1 <= ackR_unguarded(2);
      STORE_ZJ_230_store_0_ack_1 <= ackR_unguarded(1);
      STORE_ZJ_241_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_ZJ_298_word_address_0 & STORE_ZJ_230_word_address_0 & STORE_ZJ_241_word_address_0;
      data_in <= STORE_ZJ_298_data_0 & STORE_ZJ_230_data_0 & STORE_ZJ_241_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 12,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(0 downto 0),
          mdata => memory_space_1_sr_data(11 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 3,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- logger for split-operator call_stmt_275_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_275_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:call_stmt_275_call:started:  Call to module accessMem inputs: " & " konst_271_wire_constant = "& Convert_SLV_To_Hex_String(konst_271_wire_constant) & " addr_267 = "& Convert_SLV_To_Hex_String(addr_267) & " wdata_236_delayed_4_0_270 = "& Convert_SLV_To_Hex_String(wdata_236_delayed_4_0_270));
          --
        end if; 
        if call_stmt_275_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:call_stmt_275_call:finished:  outputs: " & " rdata_275= "  & Convert_SLV_To_Hex_String(rdata_275));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_330_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_330_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:call_stmt_330_call:started:  Call to module accessMem inputs: " & " konst_326_wire_constant = "& Convert_SLV_To_Hex_String(konst_326_wire_constant) & " addr_322 = "& Convert_SLV_To_Hex_String(addr_322) & " wdata_285_delayed_4_0_325 = "& Convert_SLV_To_Hex_String(wdata_285_delayed_4_0_325));
          --
        end if; 
        if call_stmt_330_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initial:DP:call_stmt_330_call:finished:  outputs: " & " rdata_330= "  & Convert_SLV_To_Hex_String(rdata_330));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_275_call call_stmt_330_call 
    accessMem_call_group_0: Block -- 
      signal data_in: std_logic_vector(57 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 10, 1 => 10);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_275_call_req_0;
      reqL_unguarded(0) <= call_stmt_330_call_req_0;
      call_stmt_275_call_ack_0 <= ackL_unguarded(1);
      call_stmt_330_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_275_call_req_1;
      reqR_unguarded(0) <= call_stmt_330_call_req_1;
      call_stmt_275_call_ack_1 <= ackR_unguarded(1);
      call_stmt_330_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessMem_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMem_call_group_0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMem_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMem_call_group_0_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMem_call_group_0_gI: SplitGuardInterface generic map(name => "accessMem_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_271_wire_constant & addr_267 & wdata_236_delayed_4_0_270 & konst_326_wire_constant & addr_322 & wdata_285_delayed_4_0_325;
      rdata_275 <= data_out(127 downto 64);
      rdata_330 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 58,
        owidth => 29,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMem_call_reqs(0),
          ackR => accessMem_call_acks(0),
          dataR => accessMem_call_data(28 downto 0),
          tagR => accessMem_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMem_return_acks(0), -- cross-over
          ackL => accessMem_return_reqs(0), -- cross-over
          dataL => accessMem_return_data(63 downto 0),
          tagL => accessMem_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end initial_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity try is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_data : out  std_logic_vector(3 downto 0);
    memory_space_8_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sc_tag :  in  std_logic_vector(0 downto 0);
    start_pipe_read_req : out  std_logic_vector(0 downto 0);
    start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    start_pipe_read_data : in   std_logic_vector(15 downto 0);
    status_pipe_write_req : out  std_logic_vector(0 downto 0);
    status_pipe_write_ack : in   std_logic_vector(0 downto 0);
    status_pipe_write_data : out  std_logic_vector(15 downto 0);
    accessMem_call_reqs : out  std_logic_vector(1 downto 0);
    accessMem_call_acks : in   std_logic_vector(1 downto 0);
    accessMem_call_data : out  std_logic_vector(57 downto 0);
    accessMem_call_tag  :  out  std_logic_vector(3 downto 0);
    accessMem_return_reqs : out  std_logic_vector(1 downto 0);
    accessMem_return_acks : in   std_logic_vector(1 downto 0);
    accessMem_return_data : in   std_logic_vector(127 downto 0);
    accessMem_return_tag :  in   std_logic_vector(3 downto 0);
    initial_call_reqs : out  std_logic_vector(0 downto 0);
    initial_call_acks : in   std_logic_vector(0 downto 0);
    initial_call_tag  :  out  std_logic_vector(0 downto 0);
    initial_return_reqs : out  std_logic_vector(0 downto 0);
    initial_return_acks : in   std_logic_vector(0 downto 0);
    initial_return_tag :  in   std_logic_vector(0 downto 0);
    try1_call_reqs : out  std_logic_vector(0 downto 0);
    try1_call_acks : in   std_logic_vector(0 downto 0);
    try1_call_tag  :  out  std_logic_vector(0 downto 0);
    try1_return_reqs : out  std_logic_vector(0 downto 0);
    try1_return_acks : in   std_logic_vector(0 downto 0);
    try1_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity try;
architecture try_arch of try is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal try_CP_4898_start: Boolean;
  signal try_CP_4898_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(11 downto 0);
      write_data : in  std_logic_vector(15 downto 0);
      read_datal : out  std_logic_vector(63 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component initial is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(11 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(11 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      accessMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessMem_call_acks : in   std_logic_vector(0 downto 0);
      accessMem_call_data : out  std_logic_vector(28 downto 0);
      accessMem_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessMem_return_acks : in   std_logic_vector(0 downto 0);
      accessMem_return_data : in   std_logic_vector(63 downto 0);
      accessMem_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component try1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(11 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(3 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(1 downto 0);
      acc_mem_pipe_write_req : out  std_logic_vector(0 downto 0);
      acc_mem_pipe_write_ack : in   std_logic_vector(0 downto 0);
      acc_mem_pipe_write_data : out  std_logic_vector(15 downto 0);
      acc_mem_add_pipe_write_req : out  std_logic_vector(0 downto 0);
      acc_mem_add_pipe_write_ack : in   std_logic_vector(0 downto 0);
      acc_mem_add_pipe_write_data : out  std_logic_vector(15 downto 0);
      accessMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessMem_call_acks : in   std_logic_vector(0 downto 0);
      accessMem_call_data : out  std_logic_vector(28 downto 0);
      accessMem_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessMem_return_acks : in   std_logic_vector(0 downto 0);
      accessMem_return_data : in   std_logic_vector(63 downto 0);
      accessMem_return_tag :  in   std_logic_vector(1 downto 0);
      accessMem_v_call_reqs : out  std_logic_vector(0 downto 0);
      accessMem_v_call_acks : in   std_logic_vector(0 downto 0);
      accessMem_v_call_data : out  std_logic_vector(28 downto 0);
      accessMem_v_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMem_v_return_reqs : out  std_logic_vector(0 downto 0);
      accessMem_v_return_acks : in   std_logic_vector(0 downto 0);
      accessMem_v_return_data : in   std_logic_vector(63 downto 0);
      accessMem_v_return_tag :  in   std_logic_vector(0 downto 0);
      accMemAccessDaemon_call_reqs : out  std_logic_vector(0 downto 0);
      accMemAccessDaemon_call_acks : in   std_logic_vector(0 downto 0);
      accMemAccessDaemon_call_data : out  std_logic_vector(31 downto 0);
      accMemAccessDaemon_call_tag  :  out  std_logic_vector(1 downto 0);
      accMemAccessDaemon_return_reqs : out  std_logic_vector(0 downto 0);
      accMemAccessDaemon_return_acks : in   std_logic_vector(0 downto 0);
      accMemAccessDaemon_return_data : in   std_logic_vector(63 downto 0);
      accMemAccessDaemon_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_758_call_req_0 : boolean;
  signal RPIPE_start_760_inst_req_0 : boolean;
  signal call_stmt_758_call_ack_1 : boolean;
  signal call_stmt_758_call_ack_0 : boolean;
  signal STORE_one_755_store_0_ack_1 : boolean;
  signal call_stmt_758_call_req_1 : boolean;
  signal STORE_zer_752_store_0_ack_1 : boolean;
  signal STORE_one_755_store_0_ack_0 : boolean;
  signal STORE_zer_752_store_0_ack_0 : boolean;
  signal STORE_zer_752_store_0_req_0 : boolean;
  signal STORE_zer_752_store_0_req_1 : boolean;
  signal NC_804_774_buf_req_1 : boolean;
  signal NC_804_774_buf_ack_1 : boolean;
  signal STORE_one_755_store_0_req_1 : boolean;
  signal phi_stmt_770_req_0 : boolean;
  signal RPIPE_start_760_inst_req_1 : boolean;
  signal phi_stmt_770_ack_0 : boolean;
  signal RPIPE_start_760_inst_ack_1 : boolean;
  signal WPIPE_status_776_inst_req_0 : boolean;
  signal WPIPE_status_776_inst_ack_0 : boolean;
  signal phi_stmt_770_req_1 : boolean;
  signal call_stmt_779_call_req_0 : boolean;
  signal call_stmt_779_call_ack_0 : boolean;
  signal NC_804_774_buf_req_0 : boolean;
  signal NC_804_774_buf_ack_0 : boolean;
  signal RPIPE_start_760_inst_ack_0 : boolean;
  signal call_stmt_766_call_req_1 : boolean;
  signal call_stmt_766_call_ack_1 : boolean;
  signal STORE_one_755_store_0_req_0 : boolean;
  signal do_while_stmt_768_branch_req_0 : boolean;
  signal call_stmt_766_call_req_0 : boolean;
  signal call_stmt_766_call_ack_0 : boolean;
  signal call_stmt_779_call_req_1 : boolean;
  signal call_stmt_779_call_ack_1 : boolean;
  signal WPIPE_status_780_inst_req_0 : boolean;
  signal WPIPE_status_780_inst_ack_0 : boolean;
  signal WPIPE_status_780_inst_req_1 : boolean;
  signal WPIPE_status_780_inst_ack_1 : boolean;
  signal WPIPE_status_776_inst_req_1 : boolean;
  signal WPIPE_status_776_inst_ack_1 : boolean;
  signal call_stmt_787_call_req_0 : boolean;
  signal call_stmt_787_call_ack_0 : boolean;
  signal call_stmt_787_call_req_1 : boolean;
  signal call_stmt_787_call_ack_1 : boolean;
  signal slice_790_inst_req_0 : boolean;
  signal slice_790_inst_ack_0 : boolean;
  signal slice_790_inst_req_1 : boolean;
  signal slice_790_inst_ack_1 : boolean;
  signal SUB_u16_u16_795_inst_req_0 : boolean;
  signal SUB_u16_u16_795_inst_ack_0 : boolean;
  signal SUB_u16_u16_795_inst_req_1 : boolean;
  signal SUB_u16_u16_795_inst_ack_1 : boolean;
  signal call_stmt_801_call_req_0 : boolean;
  signal call_stmt_801_call_ack_0 : boolean;
  signal call_stmt_801_call_req_1 : boolean;
  signal call_stmt_801_call_ack_1 : boolean;
  signal W_NC_802_inst_req_0 : boolean;
  signal W_NC_802_inst_ack_0 : boolean;
  signal W_NC_802_inst_req_1 : boolean;
  signal W_NC_802_inst_ack_1 : boolean;
  signal do_while_stmt_768_branch_ack_0 : boolean;
  signal do_while_stmt_768_branch_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "try_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  try_CP_4898_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "try_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= try_CP_4898_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= try_CP_4898_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= try_CP_4898_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,try_CP_4898_start,"try cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,try_CP_4898_symbol, "try cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  try_CP_4898: Block -- control-path 
    signal try_CP_4898_elements: BooleanArray(77 downto 0);
    -- 
  begin -- 
    try_CP_4898_elements(0) <= try_CP_4898_start;
    try_CP_4898_symbol <= try_CP_4898_elements(13);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	10 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	7 
    -- CP-element group 0:  members (46) 
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/call_stmt_758_Sample/crr
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/call_stmt_766_update_start_
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_Update/$entry
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/RPIPE_start_760_Sample/rr
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_Sample/STORE_zer_752_Split/split_ack
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_Sample/STORE_zer_752_Split/split_req
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/call_stmt_758_Update/$entry
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_Sample/STORE_zer_752_Split/$exit
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/RPIPE_start_760_sample_start_
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_Sample/STORE_zer_752_Split/$entry
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/RPIPE_start_760_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/call_stmt_758_Update/ccr
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/call_stmt_758_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_update_start_
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_sample_start_
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/$entry
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_update_start_
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_Sample/STORE_one_755_Split/split_req
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_sample_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/call_stmt_758_update_start_
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/call_stmt_758_sample_start_
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_Sample/STORE_one_755_Split/$entry
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_Update/$entry
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/call_stmt_766_Update/$entry
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/call_stmt_766_Update/ccr
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_Sample/STORE_one_755_Split/$exit
      -- CP-element group 0: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_Sample/STORE_one_755_Split/split_ack
      -- 
    -- logger for CP element group try_CP_4898_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:STORE_zer_752_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:STORE_zer_752_store_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:STORE_one_755_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:STORE_one_755_store_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:call_stmt_758_call_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:call_stmt_758_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:RPIPE_start_760_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:call_stmt_766_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_4935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(0), ack => STORE_zer_752_store_0_req_1); -- 
    rr_4924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(0), ack => STORE_zer_752_store_0_req_0); -- 
    cr_4968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(0), ack => STORE_one_755_store_0_req_1); -- 
    rr_4957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(0), ack => STORE_one_755_store_0_req_0); -- 
    crr_4977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(0), ack => call_stmt_758_call_req_0); -- 
    ccr_4982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(0), ack => call_stmt_758_call_req_1); -- 
    rr_4991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(0), ack => RPIPE_start_760_inst_req_0); -- 
    ccr_5010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(0), ack => call_stmt_766_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_Sample/word_access_start/word_0/ra
      -- CP-element group 1: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_sample_completed_
      -- 
    -- logger for CP element group try_CP_4898_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:STORE_zer_752_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_zer_752_store_0_ack_0, ack => try_CP_4898_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	12 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_update_completed_
      -- CP-element group 2: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_754_to_call_stmt_766/STORE_zer_752_Update/$exit
      -- 
    -- logger for CP element group try_CP_4898_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:STORE_zer_752_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_zer_752_store_0_ack_1, ack => try_CP_4898_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_sample_completed_
      -- CP-element group 3: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_Sample/word_access_start/word_0/ra
      -- CP-element group 3: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_Sample/word_access_start/$exit
      -- CP-element group 3: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_Sample/$exit
      -- 
    -- logger for CP element group try_CP_4898_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:STORE_one_755_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_one_755_store_0_ack_0, ack => try_CP_4898_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	12 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_Update/$exit
      -- CP-element group 4: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_Update/word_access_complete/$exit
      -- CP-element group 4: 	 assign_stmt_754_to_call_stmt_766/STORE_one_755_update_completed_
      -- 
    -- logger for CP element group try_CP_4898_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:STORE_one_755_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_one_755_store_0_ack_1, ack => try_CP_4898_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_754_to_call_stmt_766/call_stmt_758_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_754_to_call_stmt_766/call_stmt_758_Sample/cra
      -- CP-element group 5: 	 assign_stmt_754_to_call_stmt_766/call_stmt_758_sample_completed_
      -- 
    -- logger for CP element group try_CP_4898_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:call_stmt_758_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_4978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_758_call_ack_0, ack => try_CP_4898_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	11 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_754_to_call_stmt_766/call_stmt_758_update_completed_
      -- CP-element group 6: 	 assign_stmt_754_to_call_stmt_766/call_stmt_758_Update/cca
      -- CP-element group 6: 	 assign_stmt_754_to_call_stmt_766/call_stmt_758_Update/$exit
      -- 
    -- logger for CP element group try_CP_4898_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:call_stmt_758_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_4983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_758_call_ack_1, ack => try_CP_4898_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 assign_stmt_754_to_call_stmt_766/RPIPE_start_760_Update/$entry
      -- CP-element group 7: 	 assign_stmt_754_to_call_stmt_766/RPIPE_start_760_Sample/$exit
      -- CP-element group 7: 	 assign_stmt_754_to_call_stmt_766/RPIPE_start_760_update_start_
      -- CP-element group 7: 	 assign_stmt_754_to_call_stmt_766/RPIPE_start_760_sample_completed_
      -- CP-element group 7: 	 assign_stmt_754_to_call_stmt_766/RPIPE_start_760_Update/cr
      -- CP-element group 7: 	 assign_stmt_754_to_call_stmt_766/RPIPE_start_760_Sample/ra
      -- 
    -- logger for CP element group try_CP_4898_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:RPIPE_start_760_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:RPIPE_start_760_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_4992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_start_760_inst_ack_0, ack => try_CP_4898_elements(7)); -- 
    cr_4996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(7), ack => RPIPE_start_760_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	12 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_754_to_call_stmt_766/RPIPE_start_760_Update/$exit
      -- CP-element group 8: 	 assign_stmt_754_to_call_stmt_766/RPIPE_start_760_update_completed_
      -- CP-element group 8: 	 assign_stmt_754_to_call_stmt_766/RPIPE_start_760_Update/ca
      -- 
    -- logger for CP element group try_CP_4898_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:RPIPE_start_760_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_start_760_inst_ack_1, ack => try_CP_4898_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_754_to_call_stmt_766/call_stmt_766_sample_completed_
      -- CP-element group 9: 	 assign_stmt_754_to_call_stmt_766/call_stmt_766_Sample/cra
      -- CP-element group 9: 	 assign_stmt_754_to_call_stmt_766/call_stmt_766_Sample/$exit
      -- 
    -- logger for CP element group try_CP_4898_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(9) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:call_stmt_766_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_5006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_766_call_ack_0, ack => try_CP_4898_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_754_to_call_stmt_766/call_stmt_766_update_completed_
      -- CP-element group 10: 	 assign_stmt_754_to_call_stmt_766/call_stmt_766_Update/$exit
      -- CP-element group 10: 	 assign_stmt_754_to_call_stmt_766/call_stmt_766_Update/cca
      -- 
    -- logger for CP element group try_CP_4898_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:call_stmt_766_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_5011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_766_call_ack_1, ack => try_CP_4898_elements(10)); -- 
    -- CP-element group 11:  transition  output  delay-element  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	6 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (4) 
      -- CP-element group 11: 	 assign_stmt_754_to_call_stmt_766/call_stmt_766_Sample/$entry
      -- CP-element group 11: 	 assign_stmt_754_to_call_stmt_766/call_stmt_758_call_stmt_766_delay
      -- CP-element group 11: 	 assign_stmt_754_to_call_stmt_766/call_stmt_766_Sample/crr
      -- CP-element group 11: 	 assign_stmt_754_to_call_stmt_766/call_stmt_766_sample_start_
      -- 
    -- logger for CP element group try_CP_4898_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:call_stmt_766_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_5005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(11), ack => call_stmt_766_call_req_0); -- 
    -- Element group try_CP_4898_elements(11) is a control-delay.
    cp_element_11_delay: control_delay_element  generic map(name => " 11_delay", delay_value => 1)  port map(req => try_CP_4898_elements(6), ack => try_CP_4898_elements(11), clk => clk, reset =>reset);
    -- CP-element group 12:  join  transition  place  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: 	2 
    -- CP-element group 12: 	4 
    -- CP-element group 12: 	8 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 assign_stmt_754_to_call_stmt_766/$exit
      -- CP-element group 12: 	 branch_block_stmt_767/branch_block_stmt_767__entry__
      -- CP-element group 12: 	 branch_block_stmt_767/do_while_stmt_768__entry__
      -- CP-element group 12: 	 branch_block_stmt_767/$entry
      -- 
    -- logger for CP element group try_CP_4898_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    try_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= try_CP_4898_elements(10) & try_CP_4898_elements(2) & try_CP_4898_elements(4) & try_CP_4898_elements(8);
      gj_try_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_4898_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  place  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	77 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (4) 
      -- CP-element group 13: 	 $exit
      -- CP-element group 13: 	 branch_block_stmt_767/do_while_stmt_768__exit__
      -- CP-element group 13: 	 branch_block_stmt_767/$exit
      -- CP-element group 13: 	 branch_block_stmt_767/branch_block_stmt_767__exit__
      -- 
    -- logger for CP element group try_CP_4898_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    try_CP_4898_elements(13) <= try_CP_4898_elements(77);
    -- CP-element group 14:  transition  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	20 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768__entry__
      -- CP-element group 14: 	 branch_block_stmt_767/do_while_stmt_768/$entry
      -- 
    -- logger for CP element group try_CP_4898_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    try_CP_4898_elements(14) <= try_CP_4898_elements(12);
    -- CP-element group 15:  merge  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	77 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768__exit__
      -- 
    -- logger for CP element group try_CP_4898_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(15) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try_CP_4898_elements(15) is bound as output of CP function.
    -- CP-element group 16:  merge  place  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	19 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_767/do_while_stmt_768/loop_back
      -- 
    -- logger for CP element group try_CP_4898_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(16) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try_CP_4898_elements(16) is bound as output of CP function.
    -- CP-element group 17:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	22 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	75 
    -- CP-element group 17: 	76 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_767/do_while_stmt_768/condition_done
      -- CP-element group 17: 	 branch_block_stmt_767/do_while_stmt_768/loop_exit/$entry
      -- CP-element group 17: 	 branch_block_stmt_767/do_while_stmt_768/loop_taken/$entry
      -- 
    -- logger for CP element group try_CP_4898_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(17) fired."); 
        -- 
      end if; --
    end process; 
    try_CP_4898_elements(17) <= try_CP_4898_elements(22);
    -- CP-element group 18:  branch  place  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	74 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_767/do_while_stmt_768/loop_body_done
      -- 
    -- logger for CP element group try_CP_4898_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(18) fired."); 
        -- 
      end if; --
    end process; 
    try_CP_4898_elements(18) <= try_CP_4898_elements(74);
    -- CP-element group 19:  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	16 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	28 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group try_CP_4898_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(19) fired."); 
        -- 
      end if; --
    end process; 
    try_CP_4898_elements(19) <= try_CP_4898_elements(16);
    -- CP-element group 20:  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	30 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group try_CP_4898_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(20) fired."); 
        -- 
      end if; --
    end process; 
    try_CP_4898_elements(20) <= try_CP_4898_elements(14);
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	41 
    -- CP-element group 21: 	44 
    -- CP-element group 21: 	24 
    -- CP-element group 21: 	25 
    -- CP-element group 21: 	71 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/loop_body_start
      -- CP-element group 21: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/$entry
      -- 
    -- logger for CP element group try_CP_4898_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(21) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try_CP_4898_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	27 
    -- CP-element group 22: 	70 
    -- CP-element group 22: 	71 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	17 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/condition_evaluated
      -- 
    -- logger for CP element group try_CP_4898_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:do_while_stmt_768_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_5034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_5034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(22), ack => do_while_stmt_768_branch_req_0); -- 
    try_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try_CP_4898_elements(27) & try_CP_4898_elements(70) & try_CP_4898_elements(71);
      gj_try_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_4898_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	27 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/phi_stmt_770_sample_start__ps
      -- CP-element group 23: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/aggregated_phi_sample_req
      -- 
    -- logger for CP element group try_CP_4898_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(23) fired."); 
        -- 
      end if; --
    end process; 
    try_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try_CP_4898_elements(24) & try_CP_4898_elements(27);
      gj_try_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_4898_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: 	70 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	23 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/phi_stmt_770_sample_start_
      -- 
    -- logger for CP element group try_CP_4898_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(24) fired."); 
        -- 
      end if; --
    end process; 
    try_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try_CP_4898_elements(21) & try_CP_4898_elements(26) & try_CP_4898_elements(70);
      gj_try_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_4898_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	21 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	27 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/aggregated_phi_update_req
      -- CP-element group 25: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/phi_stmt_770_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/phi_stmt_770_update_start_
      -- 
    -- logger for CP element group try_CP_4898_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(25) fired."); 
        -- 
      end if; --
    end process; 
    try_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try_CP_4898_elements(21) & try_CP_4898_elements(27);
      gj_try_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_4898_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	68 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/aggregated_phi_sample_ack
      -- CP-element group 26: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/phi_stmt_770_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/phi_stmt_770_sample_completed_
      -- 
    -- logger for CP element group try_CP_4898_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(26) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try_CP_4898_elements(26) is bound as output of CP function.
    -- CP-element group 27:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	22 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	23 
    -- CP-element group 27: 	25 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/phi_stmt_770_update_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/phi_stmt_770_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/aggregated_phi_update_ack
      -- 
    -- logger for CP element group try_CP_4898_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(27) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try_CP_4898_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	19 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/phi_stmt_770_loopback_trigger
      -- 
    -- logger for CP element group try_CP_4898_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(28) fired."); 
        -- 
      end if; --
    end process; 
    try_CP_4898_elements(28) <= try_CP_4898_elements(19);
    -- CP-element group 29:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/phi_stmt_770_loopback_sample_req
      -- CP-element group 29: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/phi_stmt_770_loopback_sample_req_ps
      -- 
    -- logger for CP element group try_CP_4898_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:phi_stmt_770_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_770_loopback_sample_req_5049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_770_loopback_sample_req_5049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(29), ack => phi_stmt_770_req_1); -- 
    -- Element group try_CP_4898_elements(29) is bound as output of CP function.
    -- CP-element group 30:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	20 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/phi_stmt_770_entry_trigger
      -- 
    -- logger for CP element group try_CP_4898_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(30) fired."); 
        -- 
      end if; --
    end process; 
    try_CP_4898_elements(30) <= try_CP_4898_elements(20);
    -- CP-element group 31:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/phi_stmt_770_entry_sample_req
      -- CP-element group 31: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/phi_stmt_770_entry_sample_req_ps
      -- 
    -- logger for CP element group try_CP_4898_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:phi_stmt_770_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_770_entry_sample_req_5052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_770_entry_sample_req_5052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(31), ack => phi_stmt_770_req_0); -- 
    -- Element group try_CP_4898_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/phi_stmt_770_phi_mux_ack
      -- CP-element group 32: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/phi_stmt_770_phi_mux_ack_ps
      -- 
    -- logger for CP element group try_CP_4898_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:phi_stmt_770_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_770_phi_mux_ack_5055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_770_ack_0, ack => try_CP_4898_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/type_cast_773_sample_start__ps
      -- CP-element group 33: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/type_cast_773_sample_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/type_cast_773_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/type_cast_773_sample_completed_
      -- 
    -- logger for CP element group try_CP_4898_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(33) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try_CP_4898_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/type_cast_773_update_start__ps
      -- CP-element group 34: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/type_cast_773_update_start_
      -- 
    -- logger for CP element group try_CP_4898_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(34) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try_CP_4898_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	36 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/type_cast_773_update_completed__ps
      -- 
    -- logger for CP element group try_CP_4898_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(35) fired."); 
        -- 
      end if; --
    end process; 
    try_CP_4898_elements(35) <= try_CP_4898_elements(36);
    -- CP-element group 36:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	35 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/type_cast_773_update_completed_
      -- 
    -- logger for CP element group try_CP_4898_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(36) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try_CP_4898_elements(36) is a control-delay.
    cp_element_36_delay: control_delay_element  generic map(name => " 36_delay", delay_value => 1)  port map(req => try_CP_4898_elements(34), ack => try_CP_4898_elements(36), clk => clk, reset =>reset);
    -- CP-element group 37:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/R_NC_774_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/R_NC_774_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/R_NC_774_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/R_NC_774_sample_start__ps
      -- 
    -- logger for CP element group try_CP_4898_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:NC_804_774_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_5076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(37), ack => NC_804_774_buf_req_0); -- 
    -- Element group try_CP_4898_elements(37) is bound as output of CP function.
    -- CP-element group 38:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/R_NC_774_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/R_NC_774_Update/req
      -- CP-element group 38: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/R_NC_774_update_start_
      -- CP-element group 38: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/R_NC_774_update_start__ps
      -- 
    -- logger for CP element group try_CP_4898_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(38) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:NC_804_774_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_5081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(38), ack => NC_804_774_buf_req_1); -- 
    -- Element group try_CP_4898_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/R_NC_774_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/R_NC_774_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/R_NC_774_Sample/ack
      -- CP-element group 39: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/R_NC_774_sample_completed__ps
      -- 
    -- logger for CP element group try_CP_4898_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:NC_804_774_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NC_804_774_buf_ack_0, ack => try_CP_4898_elements(39)); -- 
    -- CP-element group 40:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/R_NC_774_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/R_NC_774_Update/ack
      -- CP-element group 40: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/R_NC_774_update_completed__ps
      -- CP-element group 40: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/R_NC_774_update_completed_
      -- 
    -- logger for CP element group try_CP_4898_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(40) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:NC_804_774_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_5082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NC_804_774_buf_ack_1, ack => try_CP_4898_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	21 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	43 
    -- CP-element group 41: 	50 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_776_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_776_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_776_Sample/req
      -- 
    -- logger for CP element group try_CP_4898_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(41) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:WPIPE_status_776_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_5091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(41), ack => WPIPE_status_776_inst_req_0); -- 
    try_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try_CP_4898_elements(21) & try_CP_4898_elements(43) & try_CP_4898_elements(50);
      gj_try_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_4898_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_776_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_776_update_start_
      -- CP-element group 42: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_776_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_776_Sample/ack
      -- CP-element group 42: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_776_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_776_Update/req
      -- 
    -- logger for CP element group try_CP_4898_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(42) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:WPIPE_status_776_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:WPIPE_status_776_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_5092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_status_776_inst_ack_0, ack => try_CP_4898_elements(42)); -- 
    req_5096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(42), ack => WPIPE_status_776_inst_req_1); -- 
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	48 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	41 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_776_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_776_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_776_Update/ack
      -- 
    -- logger for CP element group try_CP_4898_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(43) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:WPIPE_status_776_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_5097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_status_776_inst_ack_1, ack => try_CP_4898_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	21 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	46 
    -- CP-element group 44: 	66 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_779_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_779_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_779_Sample/crr
      -- 
    -- logger for CP element group try_CP_4898_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(44) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:call_stmt_779_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_5105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(44), ack => call_stmt_779_call_req_0); -- 
    try_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 23) := "try_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try_CP_4898_elements(21) & try_CP_4898_elements(46) & try_CP_4898_elements(66);
      gj_try_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_4898_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: marked-predecessors 
    -- CP-element group 45: 	47 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_779_update_start_
      -- CP-element group 45: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_779_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_779_Update/ccr
      -- 
    -- logger for CP element group try_CP_4898_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(45) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:call_stmt_779_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_5110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(45), ack => call_stmt_779_call_req_1); -- 
    try_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try_CP_4898_elements(47);
      gj_try_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_4898_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	44 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_779_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_779_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_779_Sample/cra
      -- 
    -- logger for CP element group try_CP_4898_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(46) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:call_stmt_779_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_5106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_779_call_ack_0, ack => try_CP_4898_elements(46)); -- 
    -- CP-element group 47:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	72 
    -- CP-element group 47: marked-successors 
    -- CP-element group 47: 	45 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_779_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_779_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_779_Update/cca
      -- 
    -- logger for CP element group try_CP_4898_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(47) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:call_stmt_779_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_5111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_779_call_ack_1, ack => try_CP_4898_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	43 
    -- CP-element group 48: marked-predecessors 
    -- CP-element group 48: 	50 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_780_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_780_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_780_Sample/req
      -- 
    -- logger for CP element group try_CP_4898_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(48) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:WPIPE_status_780_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_5119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(48), ack => WPIPE_status_780_inst_req_0); -- 
    try_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try_CP_4898_elements(43) & try_CP_4898_elements(50);
      gj_try_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_4898_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_780_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_780_update_start_
      -- CP-element group 49: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_780_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_780_Sample/ack
      -- CP-element group 49: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_780_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_780_Update/req
      -- 
    -- logger for CP element group try_CP_4898_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(49) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:WPIPE_status_780_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:WPIPE_status_780_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_5120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_status_780_inst_ack_0, ack => try_CP_4898_elements(49)); -- 
    req_5124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(49), ack => WPIPE_status_780_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	74 
    -- CP-element group 50: marked-successors 
    -- CP-element group 50: 	41 
    -- CP-element group 50: 	48 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_780_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_780_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/WPIPE_status_780_Update/ack
      -- 
    -- logger for CP element group try_CP_4898_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(50) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:WPIPE_status_780_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_5125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_status_780_inst_ack_1, ack => try_CP_4898_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	72 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	53 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_787_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_787_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_787_Sample/crr
      -- 
    -- logger for CP element group try_CP_4898_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(51) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:call_stmt_787_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_5133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(51), ack => call_stmt_787_call_req_0); -- 
    try_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 23) := "try_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try_CP_4898_elements(72) & try_CP_4898_elements(53);
      gj_try_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_4898_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: 	57 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_787_update_start_
      -- CP-element group 52: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_787_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_787_Update/ccr
      -- 
    -- logger for CP element group try_CP_4898_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(52) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:call_stmt_787_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_5138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(52), ack => call_stmt_787_call_req_1); -- 
    try_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try_CP_4898_elements(54) & try_CP_4898_elements(57);
      gj_try_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_4898_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: marked-successors 
    -- CP-element group 53: 	51 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_787_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_787_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_787_Sample/cra
      -- 
    -- logger for CP element group try_CP_4898_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(53) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:call_stmt_787_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_5134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_787_call_ack_0, ack => try_CP_4898_elements(53)); -- 
    -- CP-element group 54:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	73 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	52 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_787_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_787_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_787_Update/cca
      -- 
    -- logger for CP element group try_CP_4898_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(54) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:call_stmt_787_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_5139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_787_call_ack_1, ack => try_CP_4898_elements(54)); -- 
    -- CP-element group 55:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	57 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/slice_790_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/slice_790_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/slice_790_Sample/rr
      -- 
    -- logger for CP element group try_CP_4898_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(55) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:slice_790_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_5147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(55), ack => slice_790_inst_req_0); -- 
    try_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 23) := "try_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try_CP_4898_elements(54) & try_CP_4898_elements(57);
      gj_try_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_4898_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: 	61 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/slice_790_update_start_
      -- CP-element group 56: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/slice_790_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/slice_790_Update/cr
      -- 
    -- logger for CP element group try_CP_4898_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(56) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:slice_790_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_5152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(56), ack => slice_790_inst_req_1); -- 
    try_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try_CP_4898_elements(58) & try_CP_4898_elements(61);
      gj_try_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_4898_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	52 
    -- CP-element group 57: 	55 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/slice_790_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/slice_790_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/slice_790_Sample/ra
      -- 
    -- logger for CP element group try_CP_4898_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(57) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:slice_790_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_790_inst_ack_0, ack => try_CP_4898_elements(57)); -- 
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/slice_790_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/slice_790_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/slice_790_Update/ca
      -- 
    -- logger for CP element group try_CP_4898_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(58) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:slice_790_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_790_inst_ack_1, ack => try_CP_4898_elements(58)); -- 
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/SUB_u16_u16_795_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/SUB_u16_u16_795_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/SUB_u16_u16_795_Sample/rr
      -- 
    -- logger for CP element group try_CP_4898_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(59) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:SUB_u16_u16_795_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_5161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(59), ack => SUB_u16_u16_795_inst_req_0); -- 
    try_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 23) := "try_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try_CP_4898_elements(58) & try_CP_4898_elements(61);
      gj_try_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_4898_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: 	65 
    -- CP-element group 60: 	69 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/SUB_u16_u16_795_update_start_
      -- CP-element group 60: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/SUB_u16_u16_795_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/SUB_u16_u16_795_Update/cr
      -- 
    -- logger for CP element group try_CP_4898_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(60) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:SUB_u16_u16_795_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_5166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(60), ack => SUB_u16_u16_795_inst_req_1); -- 
    try_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try_CP_4898_elements(62) & try_CP_4898_elements(65) & try_CP_4898_elements(69);
      gj_try_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_4898_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	56 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/SUB_u16_u16_795_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/SUB_u16_u16_795_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/SUB_u16_u16_795_Sample/ra
      -- 
    -- logger for CP element group try_CP_4898_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(61) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:SUB_u16_u16_795_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_795_inst_ack_0, ack => try_CP_4898_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	67 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/SUB_u16_u16_795_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/SUB_u16_u16_795_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/SUB_u16_u16_795_Update/ca
      -- 
    -- logger for CP element group try_CP_4898_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(62) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:SUB_u16_u16_795_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_795_inst_ack_1, ack => try_CP_4898_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: 	73 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_801_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_801_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_801_Sample/crr
      -- 
    -- logger for CP element group try_CP_4898_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(63) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:call_stmt_801_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_5175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(63), ack => call_stmt_801_call_req_0); -- 
    try_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 23) := "try_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try_CP_4898_elements(62) & try_CP_4898_elements(73) & try_CP_4898_elements(65);
      gj_try_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_4898_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: marked-predecessors 
    -- CP-element group 64: 	66 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_801_update_start_
      -- CP-element group 64: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_801_Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_801_Update/ccr
      -- 
    -- logger for CP element group try_CP_4898_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(64) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:call_stmt_801_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_5180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(64), ack => call_stmt_801_call_req_1); -- 
    try_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try_CP_4898_elements(66);
      gj_try_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_4898_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: marked-successors 
    -- CP-element group 65: 	60 
    -- CP-element group 65: 	63 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_801_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_801_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_801_Sample/cra
      -- 
    -- logger for CP element group try_CP_4898_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(65) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:call_stmt_801_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_5176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_801_call_ack_0, ack => try_CP_4898_elements(65)); -- 
    -- CP-element group 66:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	74 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	44 
    -- CP-element group 66: 	64 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_801_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_801_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_801_Update/cca
      -- CP-element group 66: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/ring_reenable_memory_space_5
      -- 
    -- logger for CP element group try_CP_4898_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(66) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:call_stmt_801_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_5181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_801_call_ack_1, ack => try_CP_4898_elements(66)); -- 
    -- CP-element group 67:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	62 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/assign_stmt_804_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/assign_stmt_804_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/assign_stmt_804_Sample/req
      -- 
    -- logger for CP element group try_CP_4898_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(67) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:W_NC_802_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_5189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(67), ack => W_NC_802_inst_req_0); -- 
    try_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 23) := "try_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try_CP_4898_elements(62) & try_CP_4898_elements(69);
      gj_try_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_4898_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	26 
    -- CP-element group 68: marked-predecessors 
    -- CP-element group 68: 	70 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/assign_stmt_804_update_start_
      -- CP-element group 68: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/assign_stmt_804_Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/assign_stmt_804_Update/req
      -- 
    -- logger for CP element group try_CP_4898_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(68) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:W_NC_802_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_5194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_4898_elements(68), ack => W_NC_802_inst_req_1); -- 
    try_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try_CP_4898_elements(26) & try_CP_4898_elements(70);
      gj_try_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_4898_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	60 
    -- CP-element group 69: 	67 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/assign_stmt_804_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/assign_stmt_804_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/assign_stmt_804_Sample/ack
      -- 
    -- logger for CP element group try_CP_4898_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(69) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:W_NC_802_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_NC_802_inst_ack_0, ack => try_CP_4898_elements(69)); -- 
    -- CP-element group 70:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	22 
    -- CP-element group 70: marked-successors 
    -- CP-element group 70: 	24 
    -- CP-element group 70: 	68 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/assign_stmt_804_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/assign_stmt_804_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/assign_stmt_804_Update/ack
      -- 
    -- logger for CP element group try_CP_4898_elements(70)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(70)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(70) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:W_NC_802_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_5195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_NC_802_inst_ack_1, ack => try_CP_4898_elements(70)); -- 
    -- CP-element group 71:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	21 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	22 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group try_CP_4898_elements(71)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(71)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(71) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try_CP_4898_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => try_CP_4898_elements(21), ack => try_CP_4898_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	47 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	51 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_779_call_stmt_787_delay
      -- 
    -- logger for CP element group try_CP_4898_elements(72)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(72)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(72) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try_CP_4898_elements(72) is a control-delay.
    cp_element_72_delay: control_delay_element  generic map(name => " 72_delay", delay_value => 1)  port map(req => try_CP_4898_elements(47), ack => try_CP_4898_elements(72), clk => clk, reset =>reset);
    -- CP-element group 73:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	54 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	63 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/call_stmt_787_call_stmt_801_delay
      -- 
    -- logger for CP element group try_CP_4898_elements(73)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(73)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(73) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try_CP_4898_elements(73) is a control-delay.
    cp_element_73_delay: control_delay_element  generic map(name => " 73_delay", delay_value => 1)  port map(req => try_CP_4898_elements(54), ack => try_CP_4898_elements(73), clk => clk, reset =>reset);
    -- CP-element group 74:  join  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	50 
    -- CP-element group 74: 	66 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	18 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_767/do_while_stmt_768/do_while_stmt_768_loop_body/$exit
      -- 
    -- logger for CP element group try_CP_4898_elements(74)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(74)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(74) fired."); 
        -- 
      end if; --
    end process; 
    try_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try_CP_4898_elements(50) & try_CP_4898_elements(66);
      gj_try_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_4898_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	17 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_767/do_while_stmt_768/loop_exit/$exit
      -- CP-element group 75: 	 branch_block_stmt_767/do_while_stmt_768/loop_exit/ack
      -- 
    -- logger for CP element group try_CP_4898_elements(75)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(75)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(75) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:do_while_stmt_768_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_768_branch_ack_0, ack => try_CP_4898_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	17 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_767/do_while_stmt_768/loop_taken/$exit
      -- CP-element group 76: 	 branch_block_stmt_767/do_while_stmt_768/loop_taken/ack
      -- 
    -- logger for CP element group try_CP_4898_elements(76)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(76)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(76) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:do_while_stmt_768_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_5207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_768_branch_ack_1, ack => try_CP_4898_elements(76)); -- 
    -- CP-element group 77:  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	15 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	13 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_767/do_while_stmt_768/$exit
      -- 
    -- logger for CP element group try_CP_4898_elements(77)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try_CP_4898_elements(77)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try:CP:try_CP_4898_elements(77) fired."); 
        -- 
      end if; --
    end process; 
    try_CP_4898_elements(77) <= try_CP_4898_elements(15);
    try_do_while_stmt_768_terminator_5208: loop_terminator -- 
      generic map (name => " try_do_while_stmt_768_terminator_5208", max_iterations_in_flight =>7) 
      port map(loop_body_exit => try_CP_4898_elements(18),loop_continue => try_CP_4898_elements(76),loop_terminate => try_CP_4898_elements(75),loop_back => try_CP_4898_elements(16),loop_exit => try_CP_4898_elements(15),clk => clk, reset => reset); -- 
    phi_stmt_770_phi_seq_5083_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= try_CP_4898_elements(30);
      try_CP_4898_elements(33)<= src_sample_reqs(0);
      src_sample_acks(0)  <= try_CP_4898_elements(33);
      try_CP_4898_elements(34)<= src_update_reqs(0);
      src_update_acks(0)  <= try_CP_4898_elements(35);
      try_CP_4898_elements(31) <= phi_mux_reqs(0);
      triggers(1)  <= try_CP_4898_elements(28);
      try_CP_4898_elements(37)<= src_sample_reqs(1);
      src_sample_acks(1)  <= try_CP_4898_elements(39);
      try_CP_4898_elements(38)<= src_update_reqs(1);
      src_update_acks(1)  <= try_CP_4898_elements(40);
      try_CP_4898_elements(29) <= phi_mux_reqs(1);
      phi_stmt_770_phi_seq_5083 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_770_phi_seq_5083") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => try_CP_4898_elements(23), 
          phi_sample_ack => try_CP_4898_elements(26), 
          phi_update_req => try_CP_4898_elements(25), 
          phi_update_ack => try_CP_4898_elements(27), 
          phi_mux_ack => try_CP_4898_elements(32), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_5035_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= try_CP_4898_elements(19);
        preds(1)  <= try_CP_4898_elements(20);
        entry_tmerge_5035 : transition_merge -- 
          generic map(name => " entry_tmerge_5035")
          port map (preds => preds, symbol_out => try_CP_4898_elements(21));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal C_770 : std_logic_vector(15 downto 0);
    signal NC_804 : std_logic_vector(15 downto 0);
    signal NC_804_774_buffered : std_logic_vector(15 downto 0);
    signal STORE_one_755_data_0 : std_logic_vector(0 downto 0);
    signal STORE_one_755_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_zer_752_data_0 : std_logic_vector(3 downto 0);
    signal STORE_zer_752_word_address_0 : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_808_wire : std_logic_vector(0 downto 0);
    signal com0_791 : std_logic_vector(15 downto 0);
    signal konst_753_wire_constant : std_logic_vector(3 downto 0);
    signal konst_756_wire_constant : std_logic_vector(0 downto 0);
    signal konst_762_wire_constant : std_logic_vector(0 downto 0);
    signal konst_763_wire_constant : std_logic_vector(11 downto 0);
    signal konst_764_wire_constant : std_logic_vector(15 downto 0);
    signal konst_777_wire_constant : std_logic_vector(15 downto 0);
    signal konst_781_wire_constant : std_logic_vector(15 downto 0);
    signal konst_783_wire_constant : std_logic_vector(0 downto 0);
    signal konst_784_wire_constant : std_logic_vector(11 downto 0);
    signal konst_785_wire_constant : std_logic_vector(15 downto 0);
    signal konst_794_wire_constant : std_logic_vector(15 downto 0);
    signal konst_797_wire_constant : std_logic_vector(0 downto 0);
    signal konst_798_wire_constant : std_logic_vector(11 downto 0);
    signal konst_807_wire_constant : std_logic_vector(15 downto 0);
    signal rdatacom1_766 : std_logic_vector(63 downto 0);
    signal rdatacom2_801 : std_logic_vector(63 downto 0);
    signal rdatacom_787 : std_logic_vector(63 downto 0);
    signal star_761 : std_logic_vector(15 downto 0);
    signal type_cast_773_wire_constant : std_logic_vector(15 downto 0);
    signal wdatacom2_796 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    STORE_one_755_word_address_0 <= "0";
    STORE_zer_752_word_address_0 <= "0";
    konst_753_wire_constant <= "0000";
    konst_756_wire_constant <= "1";
    konst_762_wire_constant <= "0";
    konst_763_wire_constant <= "010000010000";
    konst_764_wire_constant <= "0000000000000001";
    konst_777_wire_constant <= "0000000000000000";
    konst_781_wire_constant <= "0000000000000001";
    konst_783_wire_constant <= "1";
    konst_784_wire_constant <= "010000010000";
    konst_785_wire_constant <= "0000000000000000";
    konst_794_wire_constant <= "0000000000000001";
    konst_797_wire_constant <= "0";
    konst_798_wire_constant <= "010000010000";
    konst_807_wire_constant <= "0000000000000000";
    type_cast_773_wire_constant <= "0000000000000000";
    -- logger for phi phi_stmt_770
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_770_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:try:DP:phi_stmt_770:input-0 type_cast_773_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_773_wire_constant));
          --
        end if;
        if phi_stmt_770_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:try:DP:phi_stmt_770:input-1 NC_804_774_buffered= " & Convert_SLV_To_Hex_String(NC_804_774_buffered));
          --
        end if;
        if phi_stmt_770_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:try:DP:phi_stmt_770:sample-completed");
          --
        end if;
        if phi_stmt_770_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:try:DP:phi_stmt_770:output C_770= " & Convert_SLV_To_Hex_String(C_770));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_770: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_773_wire_constant & NC_804_774_buffered;
      req <= phi_stmt_770_req_0 & phi_stmt_770_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_770",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_770_ack_0,
          idata => idata,
          odata => C_770,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_770
    -- logger for split-operator slice_790_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_790_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:slice_790_inst:started:   inputs: " & " rdatacom_787 = "& Convert_SLV_To_Hex_String(rdatacom_787));
          --
        end if; 
        if slice_790_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:slice_790_inst:finished:  outputs: " & " com0_791= "  & Convert_SLV_To_Hex_String(com0_791));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_790_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_790_inst_req_0;
      slice_790_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_790_inst_req_1;
      slice_790_inst_ack_1<= update_ack(0);
      slice_790_inst: SliceSplitProtocol generic map(name => "slice_790_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => rdatacom_787, dout => com0_791, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator NC_804_774_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if NC_804_774_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:NC_804_774_buf:started:   inputs: " & " NC_804 = "& Convert_SLV_To_Hex_String(NC_804));
          --
        end if; 
        if NC_804_774_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:NC_804_774_buf:finished:  outputs: " & " NC_804_774_buffered= "  & Convert_SLV_To_Hex_String(NC_804_774_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    NC_804_774_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= NC_804_774_buf_req_0;
      NC_804_774_buf_ack_0<= wack(0);
      rreq(0) <= NC_804_774_buf_req_1;
      NC_804_774_buf_ack_1<= rack(0);
      NC_804_774_buf : InterlockBuffer generic map ( -- 
        name => "NC_804_774_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => NC_804,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NC_804_774_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_NC_802_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_NC_802_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:W_NC_802_inst:started:   inputs: " & " wdatacom2_796 = "& Convert_SLV_To_Hex_String(wdatacom2_796));
          --
        end if; 
        if W_NC_802_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:W_NC_802_inst:finished:  outputs: " & " NC_804= "  & Convert_SLV_To_Hex_String(NC_804));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_NC_802_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_NC_802_inst_req_0;
      W_NC_802_inst_ack_0<= wack(0);
      rreq(0) <= W_NC_802_inst_req_1;
      W_NC_802_inst_ack_1<= rack(0);
      W_NC_802_inst : InterlockBuffer generic map ( -- 
        name => "W_NC_802_inst",
        buffer_size => 2,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => wdatacom2_796,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NC_804,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for operator STORE_one_755_gather_scatter flow-through 
    process(STORE_one_755_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:STORE_one_755_gather_scatter:flowthrough  inputs: " & " konst_756_wire_constant = "& Convert_SLV_To_Hex_String(konst_756_wire_constant) & "outputs: " & " STORE_one_755_data_0= "  & Convert_SLV_To_Hex_String(STORE_one_755_data_0));
      --
    end process; 
    -- equivalence STORE_one_755_gather_scatter
    process(konst_756_wire_constant) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := konst_756_wire_constant;
      ov(0 downto 0) := iv;
      STORE_one_755_data_0 <= ov(0 downto 0);
      --
    end process;
    -- logger for operator STORE_zer_752_gather_scatter flow-through 
    process(STORE_zer_752_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:STORE_zer_752_gather_scatter:flowthrough  inputs: " & " konst_753_wire_constant = "& Convert_SLV_To_Hex_String(konst_753_wire_constant) & "outputs: " & " STORE_zer_752_data_0= "  & Convert_SLV_To_Hex_String(STORE_zer_752_data_0));
      --
    end process; 
    -- equivalence STORE_zer_752_gather_scatter
    process(konst_753_wire_constant) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := konst_753_wire_constant;
      ov(3 downto 0) := iv;
      STORE_zer_752_data_0 <= ov(3 downto 0);
      --
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_768_branch_req_0," req0 do_while_stmt_768_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_768_branch_ack_0," ack0 do_while_stmt_768_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_768_branch_ack_1," ack1 do_while_stmt_768_branch");
    do_while_stmt_768_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= UGT_u16_u1_808_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_768_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_768_branch_req_0,
          ack0 => do_while_stmt_768_branch_ack_0,
          ack1 => do_while_stmt_768_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator SUB_u16_u16_795_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if SUB_u16_u16_795_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:SUB_u16_u16_795_inst:started:   inputs: " & " com0_791 = "& Convert_SLV_To_Hex_String(com0_791) & " konst_794_wire_constant = "& Convert_SLV_To_Hex_String(konst_794_wire_constant));
          --
        end if; 
        if SUB_u16_u16_795_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:SUB_u16_u16_795_inst:finished:  outputs: " & " wdatacom2_796= "  & Convert_SLV_To_Hex_String(wdatacom2_796));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (0) : SUB_u16_u16_795_inst 
    ApIntSub_group_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= com0_791;
      wdatacom2_796 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_795_inst_req_0;
      SUB_u16_u16_795_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_795_inst_req_1;
      SUB_u16_u16_795_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_0_gI: SplitGuardInterface generic map(name => "ApIntSub_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- logger for split-operator UGT_u16_u1_808_inst flow-through 
    process(UGT_u16_u1_808_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:UGT_u16_u1_808_inst:flowthrough inputs: " & " NC_804 = "& Convert_SLV_To_Hex_String(NC_804) & " konst_807_wire_constant = "& Convert_SLV_To_Hex_String(konst_807_wire_constant) & " outputs:" & " UGT_u16_u1_808_wire= "  & Convert_SLV_To_Hex_String(UGT_u16_u1_808_wire));
      --
    end process; 
    -- binary operator UGT_u16_u1_808_inst
    process(NC_804) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(NC_804, konst_807_wire_constant, tmp_var);
      UGT_u16_u1_808_wire <= tmp_var; --
    end process;
    -- logger for split-operator STORE_one_755_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if STORE_one_755_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:STORE_one_755_store_0:started:   inputs: " & " STORE_one_755_word_address_0 = "& Convert_SLV_To_Hex_String(STORE_one_755_word_address_0) & " STORE_one_755_data_0 = "& Convert_SLV_To_Hex_String(STORE_one_755_data_0));
          --
        end if; 
        if STORE_one_755_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:STORE_one_755_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      STORE_one_755_store_0_req_0,
      STORE_one_755_store_0_ack_0,
      STORE_one_755_store_0_req_1,
      STORE_one_755_store_0_ack_1,
      "STORE_one_755_store_0",
      "memory_space_6" ,
      STORE_one_755_data_0,
      STORE_one_755_word_address_0,
      "STORE_one_755_data_0",
      "STORE_one_755_word_address_0" -- 
    );
    -- shared store operator group (0) : STORE_one_755_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_one_755_store_0_req_0;
      STORE_one_755_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_one_755_store_0_req_1;
      STORE_one_755_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_one_755_word_address_0;
      data_in <= STORE_one_755_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 1,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(0 downto 0),
          mdata => memory_space_6_sr_data(0 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- logger for split-operator STORE_zer_752_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if STORE_zer_752_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:STORE_zer_752_store_0:started:   inputs: " & " STORE_zer_752_word_address_0 = "& Convert_SLV_To_Hex_String(STORE_zer_752_word_address_0) & " STORE_zer_752_data_0 = "& Convert_SLV_To_Hex_String(STORE_zer_752_data_0));
          --
        end if; 
        if STORE_zer_752_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:STORE_zer_752_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      STORE_zer_752_store_0_req_0,
      STORE_zer_752_store_0_ack_0,
      STORE_zer_752_store_0_req_1,
      STORE_zer_752_store_0_ack_1,
      "STORE_zer_752_store_0",
      "memory_space_8" ,
      STORE_zer_752_data_0,
      STORE_zer_752_word_address_0,
      "STORE_zer_752_data_0",
      "STORE_zer_752_word_address_0" -- 
    );
    -- shared store operator group (1) : STORE_zer_752_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_zer_752_store_0_req_0;
      STORE_zer_752_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_zer_752_store_0_req_1;
      STORE_zer_752_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_zer_752_word_address_0;
      data_in <= STORE_zer_752_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 1,
        data_width => 4,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_8_sr_req(0),
          mack => memory_space_8_sr_ack(0),
          maddr => memory_space_8_sr_addr(0 downto 0),
          mdata => memory_space_8_sr_data(3 downto 0),
          mtag => memory_space_8_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_8_sc_req(0),
          mack => memory_space_8_sc_ack(0),
          mtag => memory_space_8_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- logger for split-operator RPIPE_start_760_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_start_760_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:RPIPE_start_760_inst:started:   PipeRead from start inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_start_760_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:RPIPE_start_760_inst:finished:  outputs: " & " star_761= "  & Convert_SLV_To_Hex_String(star_761));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_start_760_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_start_760_inst_req_0;
      RPIPE_start_760_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_start_760_inst_req_1;
      RPIPE_start_760_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      star_761 <= data_out(15 downto 0);
      start_read_0_gI: SplitGuardInterface generic map(name => "start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      start_read_0: InputPortRevised -- 
        generic map ( name => "start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => start_pipe_read_req(0),
          oack => start_pipe_read_ack(0),
          odata => start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator WPIPE_status_776_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_status_776_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:WPIPE_status_776_inst:started:   PipeWrite to status inputs: " & " konst_777_wire_constant = "& Convert_SLV_To_Hex_String(konst_777_wire_constant));
          --
        end if; 
        if WPIPE_status_776_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:WPIPE_status_776_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator WPIPE_status_780_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_status_780_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:WPIPE_status_780_inst:started:   PipeWrite to status inputs: " & " konst_781_wire_constant = "& Convert_SLV_To_Hex_String(konst_781_wire_constant));
          --
        end if; 
        if WPIPE_status_780_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:WPIPE_status_780_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_status_776_inst WPIPE_status_780_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_status_776_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_status_780_inst_req_0;
      WPIPE_status_776_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_status_780_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_status_776_inst_req_1;
      update_req_unguarded(0) <= WPIPE_status_780_inst_req_1;
      WPIPE_status_776_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_status_780_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      data_in <= konst_777_wire_constant & konst_781_wire_constant;
      status_write_0_gI: SplitGuardInterface generic map(name => "status_write_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      status_write_0: OutputPortRevised -- 
        generic map ( name => "status", data_width => 16, num_reqs => 2, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => status_pipe_write_req(0),
          oack => status_pipe_write_ack(0),
          odata => status_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logger for split-operator call_stmt_758_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_758_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:call_stmt_758_call:started:  Call to module initial inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if call_stmt_758_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:call_stmt_758_call:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_758_call 
    initial_call_group_0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_758_call_req_0;
      call_stmt_758_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_758_call_req_1;
      call_stmt_758_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      initial_call_group_0_gI: SplitGuardInterface generic map(name => "initial_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => initial_call_reqs(0),
          ackR => initial_call_acks(0),
          tagR => initial_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => initial_return_acks(0), -- cross-over
          ackL => initial_return_reqs(0), -- cross-over
          tagL => initial_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- logger for split-operator call_stmt_766_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_766_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:call_stmt_766_call:started:  Call to module accessMem inputs: " & " konst_762_wire_constant = "& Convert_SLV_To_Hex_String(konst_762_wire_constant) & " konst_763_wire_constant = "& Convert_SLV_To_Hex_String(konst_763_wire_constant) & " konst_764_wire_constant = "& Convert_SLV_To_Hex_String(konst_764_wire_constant));
          --
        end if; 
        if call_stmt_766_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:call_stmt_766_call:finished:  outputs: " & " rdatacom1_766= "  & Convert_SLV_To_Hex_String(rdatacom1_766));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (1) : call_stmt_766_call 
    accessMem_call_group_1: Block -- 
      signal data_in: std_logic_vector(28 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_766_call_req_0;
      call_stmt_766_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_766_call_req_1;
      call_stmt_766_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMem_call_group_1_gI: SplitGuardInterface generic map(name => "accessMem_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_762_wire_constant & konst_763_wire_constant & konst_764_wire_constant;
      rdatacom1_766 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 29,
        owidth => 29,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMem_call_reqs(1),
          ackR => accessMem_call_acks(1),
          dataR => accessMem_call_data(57 downto 29),
          tagR => accessMem_call_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMem_return_acks(1), -- cross-over
          ackL => accessMem_return_reqs(1), -- cross-over
          dataL => accessMem_return_data(127 downto 64),
          tagL => accessMem_return_tag(3 downto 2),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- logger for split-operator call_stmt_779_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_779_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:call_stmt_779_call:started:  Call to module try1 inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if call_stmt_779_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:call_stmt_779_call:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (2) : call_stmt_779_call 
    try1_call_group_2: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_779_call_req_0;
      call_stmt_779_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_779_call_req_1;
      call_stmt_779_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      try1_call_group_2_gI: SplitGuardInterface generic map(name => "try1_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => try1_call_reqs(0),
          ackR => try1_call_acks(0),
          tagR => try1_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => try1_return_acks(0), -- cross-over
          ackL => try1_return_reqs(0), -- cross-over
          tagL => try1_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- logger for split-operator call_stmt_787_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_787_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:call_stmt_787_call:started:  Call to module accessMem inputs: " & " konst_783_wire_constant = "& Convert_SLV_To_Hex_String(konst_783_wire_constant) & " konst_784_wire_constant = "& Convert_SLV_To_Hex_String(konst_784_wire_constant) & " konst_785_wire_constant = "& Convert_SLV_To_Hex_String(konst_785_wire_constant));
          --
        end if; 
        if call_stmt_787_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:call_stmt_787_call:finished:  outputs: " & " rdatacom_787= "  & Convert_SLV_To_Hex_String(rdatacom_787));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_801_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_801_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:call_stmt_801_call:started:  Call to module accessMem inputs: " & " konst_797_wire_constant = "& Convert_SLV_To_Hex_String(konst_797_wire_constant) & " konst_798_wire_constant = "& Convert_SLV_To_Hex_String(konst_798_wire_constant) & " wdatacom2_796 = "& Convert_SLV_To_Hex_String(wdatacom2_796));
          --
        end if; 
        if call_stmt_801_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try:DP:call_stmt_801_call:finished:  outputs: " & " rdatacom2_801= "  & Convert_SLV_To_Hex_String(rdatacom2_801));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (3) : call_stmt_787_call call_stmt_801_call 
    accessMem_call_group_3: Block -- 
      signal data_in: std_logic_vector(57 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 10, 1 => 10);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_787_call_req_0;
      reqL_unguarded(0) <= call_stmt_801_call_req_0;
      call_stmt_787_call_ack_0 <= ackL_unguarded(1);
      call_stmt_801_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_787_call_req_1;
      reqR_unguarded(0) <= call_stmt_801_call_req_1;
      call_stmt_787_call_ack_1 <= ackR_unguarded(1);
      call_stmt_801_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessMem_call_group_3_accessRegulator_0: access_regulator_base generic map (name => "accessMem_call_group_3_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMem_call_group_3_accessRegulator_1: access_regulator_base generic map (name => "accessMem_call_group_3_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMem_call_group_3_gI: SplitGuardInterface generic map(name => "accessMem_call_group_3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_783_wire_constant & konst_784_wire_constant & konst_785_wire_constant & konst_797_wire_constant & konst_798_wire_constant & wdatacom2_796;
      rdatacom_787 <= data_out(127 downto 64);
      rdatacom2_801 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 58,
        owidth => 29,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMem_call_reqs(0),
          ackR => accessMem_call_acks(0),
          dataR => accessMem_call_data(28 downto 0),
          tagR => accessMem_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMem_return_acks(0), -- cross-over
          ackL => accessMem_return_reqs(0), -- cross-over
          dataL => accessMem_return_data(63 downto 0),
          tagL => accessMem_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- 
  end Block; -- data_path
  -- 
end try_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity try1 is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(3 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(3 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(11 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(3 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(10 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(3 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_7_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sc_tag :  in  std_logic_vector(1 downto 0);
    acc_mem_pipe_write_req : out  std_logic_vector(0 downto 0);
    acc_mem_pipe_write_ack : in   std_logic_vector(0 downto 0);
    acc_mem_pipe_write_data : out  std_logic_vector(15 downto 0);
    acc_mem_add_pipe_write_req : out  std_logic_vector(0 downto 0);
    acc_mem_add_pipe_write_ack : in   std_logic_vector(0 downto 0);
    acc_mem_add_pipe_write_data : out  std_logic_vector(15 downto 0);
    accessMem_call_reqs : out  std_logic_vector(0 downto 0);
    accessMem_call_acks : in   std_logic_vector(0 downto 0);
    accessMem_call_data : out  std_logic_vector(28 downto 0);
    accessMem_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMem_return_reqs : out  std_logic_vector(0 downto 0);
    accessMem_return_acks : in   std_logic_vector(0 downto 0);
    accessMem_return_data : in   std_logic_vector(63 downto 0);
    accessMem_return_tag :  in   std_logic_vector(1 downto 0);
    accessMem_v_call_reqs : out  std_logic_vector(0 downto 0);
    accessMem_v_call_acks : in   std_logic_vector(0 downto 0);
    accessMem_v_call_data : out  std_logic_vector(28 downto 0);
    accessMem_v_call_tag  :  out  std_logic_vector(0 downto 0);
    accessMem_v_return_reqs : out  std_logic_vector(0 downto 0);
    accessMem_v_return_acks : in   std_logic_vector(0 downto 0);
    accessMem_v_return_data : in   std_logic_vector(63 downto 0);
    accessMem_v_return_tag :  in   std_logic_vector(0 downto 0);
    accMemAccessDaemon_call_reqs : out  std_logic_vector(0 downto 0);
    accMemAccessDaemon_call_acks : in   std_logic_vector(0 downto 0);
    accMemAccessDaemon_call_data : out  std_logic_vector(31 downto 0);
    accMemAccessDaemon_call_tag  :  out  std_logic_vector(1 downto 0);
    accMemAccessDaemon_return_reqs : out  std_logic_vector(0 downto 0);
    accMemAccessDaemon_return_acks : in   std_logic_vector(0 downto 0);
    accMemAccessDaemon_return_data : in   std_logic_vector(63 downto 0);
    accMemAccessDaemon_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity try1;
architecture try1_arch of try1 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal try1_CP_1680_start: Boolean;
  signal try1_CP_1680_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(11 downto 0);
      write_data : in  std_logic_vector(15 downto 0);
      read_datal : out  std_logic_vector(63 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component accessMem_v is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(11 downto 0);
      write_data : in  std_logic_vector(15 downto 0);
      read_datal : out  std_logic_vector(63 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component accMemAccessDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      acc_mem_request : in  std_logic_vector(31 downto 0);
      acc_mem_responsel : out  std_logic_vector(31 downto 0);
      acc_mem_responseh : out  std_logic_vector(31 downto 0);
      accessMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessMem_call_acks : in   std_logic_vector(0 downto 0);
      accessMem_call_data : out  std_logic_vector(28 downto 0);
      accessMem_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessMem_return_acks : in   std_logic_vector(0 downto 0);
      accessMem_return_data : in   std_logic_vector(63 downto 0);
      accessMem_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal NT_437_350_buf_ack_1 : boolean;
  signal NT_437_350_buf_req_0 : boolean;
  signal W_T_310_delayed_4_0_352_inst_ack_0 : boolean;
  signal NT_437_350_buf_ack_0 : boolean;
  signal LOAD_ZJ_357_load_0_req_1 : boolean;
  signal do_while_stmt_344_branch_req_0 : boolean;
  signal array_obj_ref_430_store_0_ack_0 : boolean;
  signal phi_stmt_346_req_1 : boolean;
  signal phi_stmt_346_ack_0 : boolean;
  signal LOAD_ZJ_357_load_0_ack_1 : boolean;
  signal W_T_310_delayed_4_0_352_inst_req_1 : boolean;
  signal phi_stmt_346_req_0 : boolean;
  signal array_obj_ref_430_store_0_req_0 : boolean;
  signal W_T_310_delayed_4_0_352_inst_req_0 : boolean;
  signal ADD_u12_u12_358_inst_req_0 : boolean;
  signal W_T_310_delayed_4_0_352_inst_ack_1 : boolean;
  signal LOAD_ZJ_357_load_0_ack_0 : boolean;
  signal LOAD_ZJ_357_load_0_req_0 : boolean;
  signal NT_437_350_buf_req_1 : boolean;
  signal array_obj_ref_430_store_0_ack_1 : boolean;
  signal array_obj_ref_430_store_0_req_1 : boolean;
  signal ADD_u12_u12_358_inst_ack_0 : boolean;
  signal ADD_u16_u16_558_inst_req_0 : boolean;
  signal ADD_u12_u12_358_inst_req_1 : boolean;
  signal ADD_u12_u12_358_inst_ack_1 : boolean;
  signal type_cast_363_inst_req_0 : boolean;
  signal type_cast_363_inst_ack_0 : boolean;
  signal type_cast_363_inst_req_1 : boolean;
  signal type_cast_363_inst_ack_1 : boolean;
  signal LOAD_PJ_556_load_0_ack_1 : boolean;
  signal ADD_u16_u16_558_inst_ack_0 : boolean;
  signal LOAD_one_366_load_0_req_0 : boolean;
  signal LOAD_one_366_load_0_ack_0 : boolean;
  signal LOAD_one_366_load_0_req_1 : boolean;
  signal LOAD_one_366_load_0_ack_1 : boolean;
  signal CONCAT_u1_u32_368_inst_req_0 : boolean;
  signal CONCAT_u1_u32_368_inst_ack_0 : boolean;
  signal CONCAT_u1_u32_368_inst_req_1 : boolean;
  signal CONCAT_u1_u32_368_inst_ack_1 : boolean;
  signal STORE_PJ_555_store_0_req_0 : boolean;
  signal STORE_PJ_555_store_0_ack_0 : boolean;
  signal LOAD_PJ_556_load_0_req_0 : boolean;
  signal ADD_u16_u16_558_inst_req_1 : boolean;
  signal call_stmt_373_call_req_0 : boolean;
  signal call_stmt_373_call_ack_0 : boolean;
  signal ADD_u16_u16_558_inst_ack_1 : boolean;
  signal call_stmt_373_call_req_1 : boolean;
  signal call_stmt_373_call_ack_1 : boolean;
  signal LOAD_PJ_556_load_0_req_1 : boolean;
  signal slice_376_inst_req_0 : boolean;
  signal slice_376_inst_ack_0 : boolean;
  signal slice_376_inst_req_1 : boolean;
  signal slice_376_inst_ack_1 : boolean;
  signal ADD_u12_u12_553_inst_req_1 : boolean;
  signal ADD_u12_u12_553_inst_req_0 : boolean;
  signal slice_380_inst_req_0 : boolean;
  signal slice_380_inst_ack_0 : boolean;
  signal slice_380_inst_req_1 : boolean;
  signal slice_380_inst_ack_1 : boolean;
  signal STORE_PJ_555_store_0_req_1 : boolean;
  signal ADD_u12_u12_385_inst_req_0 : boolean;
  signal ADD_u12_u12_385_inst_ack_0 : boolean;
  signal ADD_u12_u12_385_inst_req_1 : boolean;
  signal ADD_u12_u12_385_inst_ack_1 : boolean;
  signal W_T_341_delayed_12_0_387_inst_req_0 : boolean;
  signal W_T_341_delayed_12_0_387_inst_ack_0 : boolean;
  signal W_T_341_delayed_12_0_387_inst_req_1 : boolean;
  signal W_T_341_delayed_12_0_387_inst_ack_1 : boolean;
  signal array_obj_ref_391_store_0_req_0 : boolean;
  signal array_obj_ref_391_store_0_ack_0 : boolean;
  signal array_obj_ref_391_store_0_req_1 : boolean;
  signal array_obj_ref_391_store_0_ack_1 : boolean;
  signal LOAD_PJ_556_load_0_ack_0 : boolean;
  signal ADD_u12_u12_553_inst_ack_1 : boolean;
  signal W_TT_345_delayed_11_0_394_inst_req_0 : boolean;
  signal W_TT_345_delayed_11_0_394_inst_ack_0 : boolean;
  signal W_TT_345_delayed_11_0_394_inst_req_1 : boolean;
  signal W_TT_345_delayed_11_0_394_inst_ack_1 : boolean;
  signal ADD_u12_u12_553_inst_ack_0 : boolean;
  signal array_obj_ref_398_store_0_req_0 : boolean;
  signal array_obj_ref_398_store_0_ack_0 : boolean;
  signal array_obj_ref_398_store_0_req_1 : boolean;
  signal array_obj_ref_398_store_0_ack_1 : boolean;
  signal slice_403_inst_req_0 : boolean;
  signal slice_403_inst_ack_0 : boolean;
  signal slice_403_inst_req_1 : boolean;
  signal slice_403_inst_ack_1 : boolean;
  signal slice_407_inst_req_0 : boolean;
  signal slice_407_inst_ack_0 : boolean;
  signal slice_407_inst_req_1 : boolean;
  signal slice_407_inst_ack_1 : boolean;
  signal ADD_u12_u12_412_inst_req_0 : boolean;
  signal ADD_u12_u12_412_inst_ack_0 : boolean;
  signal ADD_u12_u12_412_inst_req_1 : boolean;
  signal ADD_u12_u12_412_inst_ack_1 : boolean;
  signal ADD_u12_u12_417_inst_req_0 : boolean;
  signal ADD_u12_u12_417_inst_ack_0 : boolean;
  signal ADD_u12_u12_417_inst_req_1 : boolean;
  signal ADD_u12_u12_417_inst_ack_1 : boolean;
  signal W_TTT_367_delayed_11_0_419_inst_req_0 : boolean;
  signal W_TTT_367_delayed_11_0_419_inst_ack_0 : boolean;
  signal W_TTT_367_delayed_11_0_419_inst_req_1 : boolean;
  signal W_TTT_367_delayed_11_0_419_inst_ack_1 : boolean;
  signal array_obj_ref_423_store_0_req_0 : boolean;
  signal array_obj_ref_423_store_0_ack_0 : boolean;
  signal array_obj_ref_423_store_0_req_1 : boolean;
  signal array_obj_ref_423_store_0_ack_1 : boolean;
  signal W_TTTT_371_delayed_11_0_426_inst_req_0 : boolean;
  signal W_TTTT_371_delayed_11_0_426_inst_ack_0 : boolean;
  signal W_TTTT_371_delayed_11_0_426_inst_req_1 : boolean;
  signal W_TTTT_371_delayed_11_0_426_inst_ack_1 : boolean;
  signal ADD_u12_u12_436_inst_req_0 : boolean;
  signal ADD_u12_u12_436_inst_ack_0 : boolean;
  signal ADD_u12_u12_436_inst_req_1 : boolean;
  signal ADD_u12_u12_436_inst_ack_1 : boolean;
  signal do_while_stmt_344_branch_ack_0 : boolean;
  signal do_while_stmt_344_branch_ack_1 : boolean;
  signal STORE_PJ_451_store_0_req_0 : boolean;
  signal STORE_PJ_451_store_0_ack_0 : boolean;
  signal STORE_PJ_451_store_0_req_1 : boolean;
  signal STORE_PJ_451_store_0_ack_1 : boolean;
  signal do_while_stmt_455_branch_req_0 : boolean;
  signal phi_stmt_457_req_1 : boolean;
  signal phi_stmt_457_req_0 : boolean;
  signal phi_stmt_457_ack_0 : boolean;
  signal NJ_554_461_buf_req_0 : boolean;
  signal NJ_554_461_buf_ack_0 : boolean;
  signal NJ_554_461_buf_req_1 : boolean;
  signal NJ_554_461_buf_ack_1 : boolean;
  signal type_cast_465_inst_req_0 : boolean;
  signal type_cast_465_inst_ack_0 : boolean;
  signal type_cast_465_inst_req_1 : boolean;
  signal type_cast_465_inst_ack_1 : boolean;
  signal type_cast_469_inst_req_0 : boolean;
  signal type_cast_469_inst_ack_0 : boolean;
  signal type_cast_469_inst_req_1 : boolean;
  signal type_cast_469_inst_ack_1 : boolean;
  signal W_NJJ_415_delayed_2_0_471_inst_req_0 : boolean;
  signal W_NJJ_415_delayed_2_0_471_inst_ack_0 : boolean;
  signal W_NJJ_415_delayed_2_0_471_inst_req_1 : boolean;
  signal W_NJJ_415_delayed_2_0_471_inst_ack_1 : boolean;
  signal LOAD_one_475_load_0_req_0 : boolean;
  signal LOAD_one_475_load_0_ack_0 : boolean;
  signal LOAD_one_475_load_0_req_1 : boolean;
  signal LOAD_one_475_load_0_ack_1 : boolean;
  signal CONCAT_u1_u32_477_inst_req_0 : boolean;
  signal CONCAT_u1_u32_477_inst_ack_0 : boolean;
  signal CONCAT_u1_u32_477_inst_req_1 : boolean;
  signal CONCAT_u1_u32_477_inst_ack_1 : boolean;
  signal W_NGG_420_delayed_4_0_479_inst_req_0 : boolean;
  signal W_NGG_420_delayed_4_0_479_inst_ack_0 : boolean;
  signal W_NGG_420_delayed_4_0_479_inst_req_1 : boolean;
  signal W_NGG_420_delayed_4_0_479_inst_ack_1 : boolean;
  signal ADD_u32_u32_485_inst_req_0 : boolean;
  signal ADD_u32_u32_485_inst_ack_0 : boolean;
  signal ADD_u32_u32_485_inst_req_1 : boolean;
  signal ADD_u32_u32_485_inst_ack_1 : boolean;
  signal call_stmt_490_call_req_0 : boolean;
  signal call_stmt_490_call_ack_0 : boolean;
  signal call_stmt_490_call_req_1 : boolean;
  signal call_stmt_490_call_ack_1 : boolean;
  signal slice_493_inst_req_0 : boolean;
  signal slice_493_inst_ack_0 : boolean;
  signal slice_493_inst_req_1 : boolean;
  signal slice_493_inst_ack_1 : boolean;
  signal slice_497_inst_req_0 : boolean;
  signal slice_497_inst_ack_0 : boolean;
  signal slice_497_inst_req_1 : boolean;
  signal slice_497_inst_ack_1 : boolean;
  signal LOAD_PJ_500_load_0_req_0 : boolean;
  signal LOAD_PJ_500_load_0_ack_0 : boolean;
  signal LOAD_PJ_500_load_0_req_1 : boolean;
  signal LOAD_PJ_500_load_0_ack_1 : boolean;
  signal ADD_u16_u16_502_inst_req_0 : boolean;
  signal ADD_u16_u16_502_inst_ack_0 : boolean;
  signal ADD_u16_u16_502_inst_req_1 : boolean;
  signal ADD_u16_u16_502_inst_ack_1 : boolean;
  signal LOAD_PJ_505_load_0_req_0 : boolean;
  signal LOAD_PJ_505_load_0_ack_0 : boolean;
  signal LOAD_PJ_505_load_0_req_1 : boolean;
  signal LOAD_PJ_505_load_0_ack_1 : boolean;
  signal STORE_PJ_555_store_0_ack_1 : boolean;
  signal ADD_u12_u12_651_inst_req_1 : boolean;
  signal phi_stmt_642_req_1 : boolean;
  signal ADD_u12_u12_651_inst_ack_1 : boolean;
  signal array_obj_ref_508_store_0_req_0 : boolean;
  signal array_obj_ref_508_store_0_ack_0 : boolean;
  signal array_obj_ref_508_store_0_req_1 : boolean;
  signal array_obj_ref_508_store_0_ack_1 : boolean;
  signal phi_stmt_642_ack_0 : boolean;
  signal W_PPJ_444_delayed_6_0_511_inst_req_0 : boolean;
  signal W_PPJ_444_delayed_6_0_511_inst_ack_0 : boolean;
  signal W_PPJ_444_delayed_6_0_511_inst_req_1 : boolean;
  signal W_PPJ_444_delayed_6_0_511_inst_ack_1 : boolean;
  signal do_while_stmt_640_branch_req_0 : boolean;
  signal W_H_574_delayed_5_0_653_inst_ack_1 : boolean;
  signal array_obj_ref_515_store_0_req_0 : boolean;
  signal array_obj_ref_515_store_0_ack_0 : boolean;
  signal array_obj_ref_515_store_0_req_1 : boolean;
  signal array_obj_ref_515_store_0_ack_1 : boolean;
  signal slice_520_inst_req_0 : boolean;
  signal slice_520_inst_ack_0 : boolean;
  signal slice_520_inst_req_1 : boolean;
  signal slice_520_inst_ack_1 : boolean;
  signal slice_524_inst_req_0 : boolean;
  signal slice_524_inst_ack_0 : boolean;
  signal W_H_574_delayed_5_0_653_inst_req_0 : boolean;
  signal slice_524_inst_req_1 : boolean;
  signal slice_524_inst_ack_1 : boolean;
  signal LOAD_PJ_527_load_0_req_0 : boolean;
  signal LOAD_PJ_527_load_0_ack_0 : boolean;
  signal W_H_574_delayed_5_0_653_inst_ack_0 : boolean;
  signal LOAD_PJ_527_load_0_req_1 : boolean;
  signal LOAD_PJ_527_load_0_ack_1 : boolean;
  signal ADD_u16_u16_529_inst_req_0 : boolean;
  signal ADD_u16_u16_529_inst_ack_0 : boolean;
  signal ADD_u16_u16_529_inst_req_1 : boolean;
  signal ADD_u16_u16_529_inst_ack_1 : boolean;
  signal array_obj_ref_659_load_0_req_0 : boolean;
  signal W_H_574_delayed_5_0_653_inst_req_1 : boolean;
  signal LOAD_PJ_532_load_0_req_0 : boolean;
  signal LOAD_PJ_532_load_0_ack_0 : boolean;
  signal LOAD_PJ_532_load_0_req_1 : boolean;
  signal LOAD_PJ_532_load_0_ack_1 : boolean;
  signal ADD_u16_u16_534_inst_req_0 : boolean;
  signal ADD_u16_u16_534_inst_ack_0 : boolean;
  signal ADD_u16_u16_534_inst_req_1 : boolean;
  signal ADD_u16_u16_534_inst_ack_1 : boolean;
  signal W_PPPJ_466_delayed_6_0_536_inst_req_0 : boolean;
  signal W_PPPJ_466_delayed_6_0_536_inst_ack_0 : boolean;
  signal W_PPPJ_466_delayed_6_0_536_inst_req_1 : boolean;
  signal W_PPPJ_466_delayed_6_0_536_inst_ack_1 : boolean;
  signal array_obj_ref_540_store_0_req_0 : boolean;
  signal array_obj_ref_540_store_0_ack_0 : boolean;
  signal array_obj_ref_540_store_0_req_1 : boolean;
  signal array_obj_ref_540_store_0_ack_1 : boolean;
  signal W_PPPPJ_470_delayed_6_0_543_inst_req_0 : boolean;
  signal W_PPPPJ_470_delayed_6_0_543_inst_ack_0 : boolean;
  signal W_PPPPJ_470_delayed_6_0_543_inst_req_1 : boolean;
  signal W_PPPPJ_470_delayed_6_0_543_inst_ack_1 : boolean;
  signal array_obj_ref_547_store_0_req_0 : boolean;
  signal array_obj_ref_547_store_0_ack_0 : boolean;
  signal array_obj_ref_547_store_0_req_1 : boolean;
  signal array_obj_ref_547_store_0_ack_1 : boolean;
  signal do_while_stmt_455_branch_ack_0 : boolean;
  signal do_while_stmt_455_branch_ack_1 : boolean;
  signal STORE_total_573_store_0_req_0 : boolean;
  signal STORE_total_573_store_0_ack_0 : boolean;
  signal STORE_total_573_store_0_req_1 : boolean;
  signal STORE_total_573_store_0_ack_1 : boolean;
  signal do_while_stmt_577_branch_req_0 : boolean;
  signal phi_stmt_579_req_1 : boolean;
  signal phi_stmt_579_req_0 : boolean;
  signal phi_stmt_579_ack_0 : boolean;
  signal NK_612_583_buf_req_0 : boolean;
  signal NK_612_583_buf_ack_0 : boolean;
  signal NK_612_583_buf_req_1 : boolean;
  signal NK_612_583_buf_ack_1 : boolean;
  signal array_obj_ref_587_load_0_req_0 : boolean;
  signal array_obj_ref_587_load_0_ack_0 : boolean;
  signal array_obj_ref_587_load_0_req_1 : boolean;
  signal array_obj_ref_587_load_0_ack_1 : boolean;
  signal array_obj_ref_591_load_0_req_0 : boolean;
  signal array_obj_ref_591_load_0_ack_0 : boolean;
  signal array_obj_ref_591_load_0_req_1 : boolean;
  signal array_obj_ref_591_load_0_ack_1 : boolean;
  signal W_K_517_delayed_5_0_593_inst_req_0 : boolean;
  signal W_K_517_delayed_5_0_593_inst_ack_0 : boolean;
  signal W_K_517_delayed_5_0_593_inst_req_1 : boolean;
  signal W_K_517_delayed_5_0_593_inst_ack_1 : boolean;
  signal MUL_u16_u16_600_inst_req_0 : boolean;
  signal MUL_u16_u16_600_inst_ack_0 : boolean;
  signal MUL_u16_u16_600_inst_req_1 : boolean;
  signal MUL_u16_u16_600_inst_ack_1 : boolean;
  signal array_obj_ref_597_store_0_req_0 : boolean;
  signal array_obj_ref_597_store_0_ack_0 : boolean;
  signal array_obj_ref_597_store_0_req_1 : boolean;
  signal array_obj_ref_597_store_0_ack_1 : boolean;
  signal LOAD_total_603_load_0_req_0 : boolean;
  signal LOAD_total_603_load_0_ack_0 : boolean;
  signal ADD_u12_u12_651_inst_ack_0 : boolean;
  signal ADD_u12_u12_651_inst_req_0 : boolean;
  signal LOAD_total_603_load_0_req_1 : boolean;
  signal LOAD_total_603_load_0_ack_1 : boolean;
  signal NH_691_646_buf_ack_1 : boolean;
  signal NH_691_646_buf_req_1 : boolean;
  signal array_obj_ref_605_load_0_req_0 : boolean;
  signal array_obj_ref_605_load_0_ack_0 : boolean;
  signal NH_691_646_buf_ack_0 : boolean;
  signal NH_691_646_buf_req_0 : boolean;
  signal array_obj_ref_605_load_0_req_1 : boolean;
  signal array_obj_ref_605_load_0_ack_1 : boolean;
  signal array_obj_ref_659_load_0_req_1 : boolean;
  signal array_obj_ref_659_load_0_ack_1 : boolean;
  signal ADD_u16_u16_606_inst_req_0 : boolean;
  signal ADD_u16_u16_606_inst_ack_0 : boolean;
  signal ADD_u16_u16_606_inst_req_1 : boolean;
  signal ADD_u16_u16_606_inst_ack_1 : boolean;
  signal phi_stmt_642_req_0 : boolean;
  signal STORE_total_602_store_0_req_0 : boolean;
  signal STORE_total_602_store_0_ack_0 : boolean;
  signal STORE_total_602_store_0_req_1 : boolean;
  signal STORE_total_602_store_0_ack_1 : boolean;
  signal ADD_u32_u32_611_inst_req_0 : boolean;
  signal ADD_u32_u32_611_inst_ack_0 : boolean;
  signal ADD_u32_u32_611_inst_req_1 : boolean;
  signal ADD_u32_u32_611_inst_ack_1 : boolean;
  signal array_obj_ref_659_load_0_ack_0 : boolean;
  signal do_while_stmt_577_branch_ack_0 : boolean;
  signal do_while_stmt_577_branch_ack_1 : boolean;
  signal ADD_u12_u12_621_inst_req_0 : boolean;
  signal ADD_u12_u12_621_inst_ack_0 : boolean;
  signal ADD_u12_u12_621_inst_req_1 : boolean;
  signal ADD_u12_u12_621_inst_ack_1 : boolean;
  signal LOAD_total_622_load_0_req_0 : boolean;
  signal LOAD_total_622_load_0_ack_0 : boolean;
  signal LOAD_total_622_load_0_req_1 : boolean;
  signal LOAD_total_622_load_0_ack_1 : boolean;
  signal call_stmt_624_call_req_0 : boolean;
  signal call_stmt_624_call_ack_0 : boolean;
  signal call_stmt_624_call_req_1 : boolean;
  signal call_stmt_624_call_ack_1 : boolean;
  signal LOAD_zer_626_load_0_req_0 : boolean;
  signal LOAD_zer_626_load_0_ack_0 : boolean;
  signal LOAD_zer_626_load_0_req_1 : boolean;
  signal LOAD_zer_626_load_0_ack_1 : boolean;
  signal CONCAT_u4_u16_630_inst_req_0 : boolean;
  signal CONCAT_u4_u16_630_inst_ack_0 : boolean;
  signal CONCAT_u4_u16_630_inst_req_1 : boolean;
  signal CONCAT_u4_u16_630_inst_ack_1 : boolean;
  signal WPIPE_acc_mem_add_632_inst_req_0 : boolean;
  signal WPIPE_acc_mem_add_632_inst_ack_0 : boolean;
  signal WPIPE_acc_mem_add_632_inst_req_1 : boolean;
  signal WPIPE_acc_mem_add_632_inst_ack_1 : boolean;
  signal array_obj_ref_637_load_0_req_0 : boolean;
  signal array_obj_ref_637_load_0_ack_0 : boolean;
  signal array_obj_ref_637_load_0_req_1 : boolean;
  signal array_obj_ref_637_load_0_ack_1 : boolean;
  signal WPIPE_acc_mem_635_inst_req_0 : boolean;
  signal WPIPE_acc_mem_635_inst_ack_0 : boolean;
  signal WPIPE_acc_mem_635_inst_req_1 : boolean;
  signal WPIPE_acc_mem_635_inst_ack_1 : boolean;
  signal array_obj_ref_657_store_0_req_0 : boolean;
  signal array_obj_ref_657_store_0_ack_0 : boolean;
  signal array_obj_ref_657_store_0_req_1 : boolean;
  signal array_obj_ref_657_store_0_ack_1 : boolean;
  signal ADD_u12_u12_664_inst_req_0 : boolean;
  signal ADD_u12_u12_664_inst_ack_0 : boolean;
  signal ADD_u12_u12_664_inst_req_1 : boolean;
  signal ADD_u12_u12_664_inst_ack_1 : boolean;
  signal W_HH_584_delayed_4_0_666_inst_req_0 : boolean;
  signal W_HH_584_delayed_4_0_666_inst_ack_0 : boolean;
  signal W_HH_584_delayed_4_0_666_inst_req_1 : boolean;
  signal W_HH_584_delayed_4_0_666_inst_ack_1 : boolean;
  signal array_obj_ref_672_load_0_req_0 : boolean;
  signal array_obj_ref_672_load_0_ack_0 : boolean;
  signal array_obj_ref_672_load_0_req_1 : boolean;
  signal array_obj_ref_672_load_0_ack_1 : boolean;
  signal array_obj_ref_670_store_0_req_0 : boolean;
  signal array_obj_ref_670_store_0_ack_0 : boolean;
  signal array_obj_ref_670_store_0_req_1 : boolean;
  signal array_obj_ref_670_store_0_ack_1 : boolean;
  signal ADD_u12_u12_677_inst_req_0 : boolean;
  signal ADD_u12_u12_677_inst_ack_0 : boolean;
  signal ADD_u12_u12_677_inst_req_1 : boolean;
  signal ADD_u12_u12_677_inst_ack_1 : boolean;
  signal W_HHH_594_delayed_4_0_679_inst_req_0 : boolean;
  signal W_HHH_594_delayed_4_0_679_inst_ack_0 : boolean;
  signal W_HHH_594_delayed_4_0_679_inst_req_1 : boolean;
  signal W_HHH_594_delayed_4_0_679_inst_ack_1 : boolean;
  signal array_obj_ref_685_load_0_req_0 : boolean;
  signal array_obj_ref_685_load_0_ack_0 : boolean;
  signal array_obj_ref_685_load_0_req_1 : boolean;
  signal array_obj_ref_685_load_0_ack_1 : boolean;
  signal array_obj_ref_683_store_0_req_0 : boolean;
  signal array_obj_ref_683_store_0_ack_0 : boolean;
  signal array_obj_ref_683_store_0_req_1 : boolean;
  signal array_obj_ref_683_store_0_ack_1 : boolean;
  signal ADD_u12_u12_690_inst_req_0 : boolean;
  signal ADD_u12_u12_690_inst_ack_0 : boolean;
  signal ADD_u12_u12_690_inst_req_1 : boolean;
  signal ADD_u12_u12_690_inst_ack_1 : boolean;
  signal do_while_stmt_640_branch_ack_0 : boolean;
  signal do_while_stmt_640_branch_ack_1 : boolean;
  signal ADD_u12_u12_702_inst_req_0 : boolean;
  signal ADD_u12_u12_702_inst_ack_0 : boolean;
  signal ADD_u12_u12_702_inst_req_1 : boolean;
  signal ADD_u12_u12_702_inst_ack_1 : boolean;
  signal call_stmt_705_call_req_0 : boolean;
  signal call_stmt_705_call_ack_0 : boolean;
  signal call_stmt_705_call_req_1 : boolean;
  signal call_stmt_705_call_ack_1 : boolean;
  signal slice_709_inst_req_0 : boolean;
  signal slice_709_inst_ack_0 : boolean;
  signal slice_709_inst_req_1 : boolean;
  signal slice_709_inst_ack_1 : boolean;
  signal array_obj_ref_707_store_0_req_0 : boolean;
  signal array_obj_ref_707_store_0_ack_0 : boolean;
  signal array_obj_ref_707_store_0_req_1 : boolean;
  signal array_obj_ref_707_store_0_ack_1 : boolean;
  signal slice_714_inst_req_0 : boolean;
  signal slice_714_inst_ack_0 : boolean;
  signal slice_714_inst_req_1 : boolean;
  signal slice_714_inst_ack_1 : boolean;
  signal array_obj_ref_712_store_0_req_0 : boolean;
  signal array_obj_ref_712_store_0_ack_0 : boolean;
  signal array_obj_ref_712_store_0_req_1 : boolean;
  signal array_obj_ref_712_store_0_ack_1 : boolean;
  signal slice_719_inst_req_0 : boolean;
  signal slice_719_inst_ack_0 : boolean;
  signal slice_719_inst_req_1 : boolean;
  signal slice_719_inst_ack_1 : boolean;
  signal array_obj_ref_717_store_0_req_0 : boolean;
  signal array_obj_ref_717_store_0_ack_0 : boolean;
  signal array_obj_ref_717_store_0_req_1 : boolean;
  signal array_obj_ref_717_store_0_ack_1 : boolean;
  signal slice_724_inst_req_0 : boolean;
  signal slice_724_inst_ack_0 : boolean;
  signal slice_724_inst_req_1 : boolean;
  signal slice_724_inst_ack_1 : boolean;
  signal array_obj_ref_722_store_0_req_0 : boolean;
  signal array_obj_ref_722_store_0_ack_0 : boolean;
  signal array_obj_ref_722_store_0_req_1 : boolean;
  signal array_obj_ref_722_store_0_ack_1 : boolean;
  signal ADD_u12_u12_729_inst_req_0 : boolean;
  signal ADD_u12_u12_729_inst_ack_0 : boolean;
  signal ADD_u12_u12_729_inst_req_1 : boolean;
  signal ADD_u12_u12_729_inst_ack_1 : boolean;
  signal if_stmt_731_branch_req_0 : boolean;
  signal if_stmt_731_branch_ack_1 : boolean;
  signal if_stmt_731_branch_ack_0 : boolean;
  signal phi_stmt_567_req_0 : boolean;
  signal NL_730_571_buf_req_0 : boolean;
  signal NL_730_571_buf_ack_0 : boolean;
  signal NL_730_571_buf_req_1 : boolean;
  signal NL_730_571_buf_ack_1 : boolean;
  signal phi_stmt_567_req_1 : boolean;
  signal phi_stmt_567_ack_0 : boolean;
  signal ADD_u12_u12_741_inst_req_0 : boolean;
  signal ADD_u12_u12_741_inst_ack_0 : boolean;
  signal ADD_u12_u12_741_inst_req_1 : boolean;
  signal ADD_u12_u12_741_inst_ack_1 : boolean;
  signal if_stmt_743_branch_req_0 : boolean;
  signal if_stmt_743_branch_ack_1 : boolean;
  signal if_stmt_743_branch_ack_0 : boolean;
  signal phi_stmt_445_req_0 : boolean;
  signal NG_742_449_buf_req_0 : boolean;
  signal NG_742_449_buf_ack_0 : boolean;
  signal NG_742_449_buf_req_1 : boolean;
  signal NG_742_449_buf_ack_1 : boolean;
  signal phi_stmt_445_req_1 : boolean;
  signal phi_stmt_445_ack_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "try1_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  try1_CP_1680_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "try1_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= try1_CP_1680_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= try1_CP_1680_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= try1_CP_1680_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,try1_CP_1680_start,"try1 cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,try1_CP_1680_symbol, "try1 cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  try1_CP_1680: Block -- control-path 
    signal try1_CP_1680_elements: BooleanArray(527 downto 0);
    -- 
  begin -- 
    try1_CP_1680_elements(0) <= try1_CP_1680_start;
    try1_CP_1680_symbol <= try1_CP_1680_elements(521);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_343/$entry
      -- CP-element group 0: 	 branch_block_stmt_343/do_while_stmt_344__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_343/branch_block_stmt_343__entry__
      -- 
    -- logger for CP element group try1_CP_1680_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  branch  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	128 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	522 
    -- CP-element group 1:  members (10) 
      -- CP-element group 1: 	 branch_block_stmt_343/$exit
      -- CP-element group 1: 	 branch_block_stmt_343/branch_block_stmt_343__exit__
      -- CP-element group 1: 	 branch_block_stmt_443/branch_block_stmt_443__entry__
      -- CP-element group 1: 	 branch_block_stmt_343/do_while_stmt_344__exit__
      -- CP-element group 1: 	 branch_block_stmt_443/merge_stmt_444__entry__
      -- CP-element group 1: 	 branch_block_stmt_443/$entry
      -- CP-element group 1: 	 branch_block_stmt_443/merge_stmt_444_dead_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_443/merge_stmt_444__entry___PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_443/merge_stmt_444__entry___PhiReq/phi_stmt_445/$entry
      -- CP-element group 1: 	 branch_block_stmt_443/merge_stmt_444__entry___PhiReq/phi_stmt_445/phi_stmt_445_sources/$entry
      -- 
    -- logger for CP element group try1_CP_1680_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(1) <= try1_CP_1680_elements(128);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_343/do_while_stmt_344/$entry
      -- CP-element group 2: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344__entry__
      -- 
    -- logger for CP element group try1_CP_1680_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(2) <= try1_CP_1680_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	128 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344__exit__
      -- 
    -- logger for CP element group try1_CP_1680_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_343/do_while_stmt_344/loop_back
      -- 
    -- logger for CP element group try1_CP_1680_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	126 
    -- CP-element group 5: 	127 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_343/do_while_stmt_344/condition_done
      -- CP-element group 5: 	 branch_block_stmt_343/do_while_stmt_344/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_343/do_while_stmt_344/loop_taken/$entry
      -- 
    -- logger for CP element group try1_CP_1680_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(5) <= try1_CP_1680_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	125 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_343/do_while_stmt_344/loop_body_done
      -- 
    -- logger for CP element group try1_CP_1680_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(6) <= try1_CP_1680_elements(125);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group try1_CP_1680_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(7) <= try1_CP_1680_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group try1_CP_1680_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(8) <= try1_CP_1680_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9: 	121 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	47 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_root_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_root_address_calculated
      -- 
    -- logger for CP element group try1_CP_1680_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	120 
    -- CP-element group 10: 	121 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/condition_evaluated
      -- 
    -- logger for CP element group try1_CP_1680_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:do_while_stmt_344_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_1704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(10), ack => do_while_stmt_344_branch_req_0); -- 
    try1_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(15) & try1_CP_1680_elements(120) & try1_CP_1680_elements(121);
      gj_try1_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/phi_stmt_346_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/aggregated_phi_sample_req
      -- 
    -- logger for CP element group try1_CP_1680_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    try1_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(12) & try1_CP_1680_elements(15);
      gj_try1_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: 	120 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/phi_stmt_346_sample_start_
      -- 
    -- logger for CP element group try1_CP_1680_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    try1_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(9) & try1_CP_1680_elements(14) & try1_CP_1680_elements(120);
      gj_try1_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	119 
    -- CP-element group 13: 	95 
    -- CP-element group 13: 	99 
    -- CP-element group 13: 	31 
    -- CP-element group 13: 	67 
    -- CP-element group 13: 	71 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/phi_stmt_346_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/phi_stmt_346_update_start_
      -- CP-element group 13: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/aggregated_phi_update_req
      -- 
    -- logger for CP element group try1_CP_1680_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    try1_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= try1_CP_1680_elements(9) & try1_CP_1680_elements(119) & try1_CP_1680_elements(95) & try1_CP_1680_elements(99) & try1_CP_1680_elements(31) & try1_CP_1680_elements(67) & try1_CP_1680_elements(71);
      gj_try1_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	118 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/phi_stmt_346_sample_completed__ps
      -- CP-element group 14: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/phi_stmt_346_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/aggregated_phi_sample_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(14) is bound as output of CP function.
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: 	117 
    -- CP-element group 15: 	93 
    -- CP-element group 15: 	97 
    -- CP-element group 15: 	29 
    -- CP-element group 15: 	65 
    -- CP-element group 15: 	69 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/phi_stmt_346_update_completed__ps
      -- CP-element group 15: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/phi_stmt_346_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/aggregated_phi_update_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(15) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/phi_stmt_346_loopback_trigger
      -- 
    -- logger for CP element group try1_CP_1680_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(16) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(16) <= try1_CP_1680_elements(7);
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/phi_stmt_346_loopback_sample_req
      -- CP-element group 17: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/phi_stmt_346_loopback_sample_req_ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:phi_stmt_346_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_346_loopback_sample_req_1719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_346_loopback_sample_req_1719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(17), ack => phi_stmt_346_req_1); -- 
    -- Element group try1_CP_1680_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/phi_stmt_346_entry_trigger
      -- 
    -- logger for CP element group try1_CP_1680_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(18) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(18) <= try1_CP_1680_elements(8);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/phi_stmt_346_entry_sample_req
      -- CP-element group 19: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/phi_stmt_346_entry_sample_req_ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:phi_stmt_346_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_346_entry_sample_req_1722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_346_entry_sample_req_1722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(19), ack => phi_stmt_346_req_0); -- 
    -- Element group try1_CP_1680_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/phi_stmt_346_phi_mux_ack
      -- CP-element group 20: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/phi_stmt_346_phi_mux_ack_ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:phi_stmt_346_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_346_phi_mux_ack_1725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_346_ack_0, ack => try1_CP_1680_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/type_cast_349_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/type_cast_349_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/type_cast_349_sample_start__ps
      -- CP-element group 21: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/type_cast_349_sample_completed__ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(21) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/type_cast_349_update_start_
      -- CP-element group 22: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/type_cast_349_update_start__ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(22) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/type_cast_349_update_completed__ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(23) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(23) <= try1_CP_1680_elements(24);
    -- CP-element group 24:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	23 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/type_cast_349_update_completed_
      -- 
    -- logger for CP element group try1_CP_1680_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(24) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(24) is a control-delay.
    cp_element_24_delay: control_delay_element  generic map(name => " 24_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(22), ack => try1_CP_1680_elements(24), clk => clk, reset =>reset);
    -- CP-element group 25:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/R_NT_350_Sample/req
      -- CP-element group 25: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/R_NT_350_sample_start__ps
      -- CP-element group 25: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/R_NT_350_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/R_NT_350_Sample/$entry
      -- 
    -- logger for CP element group try1_CP_1680_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NT_437_350_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(25), ack => NT_437_350_buf_req_0); -- 
    -- Element group try1_CP_1680_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/R_NT_350_update_start__ps
      -- CP-element group 26: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/R_NT_350_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/R_NT_350_update_start_
      -- CP-element group 26: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/R_NT_350_Update/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NT_437_350_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(26), ack => NT_437_350_buf_req_1); -- 
    -- Element group try1_CP_1680_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/R_NT_350_Sample/ack
      -- CP-element group 27: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/R_NT_350_sample_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/R_NT_350_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/R_NT_350_sample_completed_
      -- 
    -- logger for CP element group try1_CP_1680_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NT_437_350_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NT_437_350_buf_ack_0, ack => try1_CP_1680_elements(27)); -- 
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/R_NT_350_Update/ack
      -- CP-element group 28: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/R_NT_350_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/R_NT_350_update_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/R_NT_350_update_completed_
      -- 
    -- logger for CP element group try1_CP_1680_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NT_437_350_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NT_437_350_buf_ack_1, ack => try1_CP_1680_elements(28)); -- 
    -- CP-element group 29:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	15 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	31 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_354_Sample/req
      -- CP-element group 29: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_354_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_354_sample_start_
      -- 
    -- logger for CP element group try1_CP_1680_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_T_310_delayed_4_0_352_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(29), ack => W_T_310_delayed_4_0_352_inst_req_0); -- 
    try1_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 24) := "try1_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(15) & try1_CP_1680_elements(31);
      gj_try1_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	39 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_354_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_354_Update/req
      -- CP-element group 30: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_354_update_start_
      -- 
    -- logger for CP element group try1_CP_1680_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_T_310_delayed_4_0_352_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(30), ack => W_T_310_delayed_4_0_352_inst_req_1); -- 
    try1_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(39);
      gj_try1_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: marked-successors 
    -- CP-element group 31: 	13 
    -- CP-element group 31: 	29 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_354_Sample/ack
      -- CP-element group 31: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_354_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_354_sample_completed_
      -- 
    -- logger for CP element group try1_CP_1680_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_T_310_delayed_4_0_352_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_T_310_delayed_4_0_352_inst_ack_0, ack => try1_CP_1680_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_354_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_354_Update/ack
      -- CP-element group 32: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_354_update_completed_
      -- 
    -- logger for CP element group try1_CP_1680_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_T_310_delayed_4_0_352_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_T_310_delayed_4_0_352_inst_ack_1, ack => try1_CP_1680_elements(32)); -- 
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: 	38 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	39 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	39 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_358_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_358_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_358_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_358_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(33), ack => ADD_u12_u12_358_inst_req_0); -- 
    try1_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 24) := "try1_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(32) & try1_CP_1680_elements(38) & try1_CP_1680_elements(39);
      gj_try1_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	43 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	40 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_358_update_start_
      -- CP-element group 34: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_358_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_358_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_358_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(34), ack => ADD_u12_u12_358_inst_req_1); -- 
    try1_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(43);
      gj_try1_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	37 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (5) 
      -- CP-element group 35: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_Sample/word_access_start/$entry
      -- CP-element group 35: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_Sample/word_access_start/word_0/$entry
      -- CP-element group 35: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_ZJ_357_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(35), ack => LOAD_ZJ_357_load_0_req_0); -- 
    try1_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 24) := "try1_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(9) & try1_CP_1680_elements(37);
      gj_try1_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	39 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_Update/word_access_complete/word_0/cr
      -- CP-element group 36: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_Update/word_access_complete/$entry
      -- CP-element group 36: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_update_start_
      -- CP-element group 36: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_Update/word_access_complete/word_0/$entry
      -- 
    -- logger for CP element group try1_CP_1680_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(36) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_ZJ_357_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(36), ack => LOAD_ZJ_357_load_0_req_1); -- 
    try1_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(39);
      gj_try1_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: marked-successors 
    -- CP-element group 37: 	35 
    -- CP-element group 37:  members (5) 
      -- CP-element group 37: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_Sample/word_access_start/$exit
      -- CP-element group 37: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_Sample/word_access_start/word_0/$exit
      -- CP-element group 37: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_ZJ_357_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ZJ_357_load_0_ack_0, ack => try1_CP_1680_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	33 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_Update/LOAD_ZJ_357_Merge/merge_ack
      -- CP-element group 38: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_Update/word_access_complete/$exit
      -- CP-element group 38: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_Update/word_access_complete/word_0/ca
      -- CP-element group 38: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_Update/LOAD_ZJ_357_Merge/$entry
      -- CP-element group 38: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_Update/LOAD_ZJ_357_Merge/$exit
      -- CP-element group 38: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_Update/LOAD_ZJ_357_Merge/merge_req
      -- CP-element group 38: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_ZJ_357_Update/word_access_complete/word_0/$exit
      -- 
    -- logger for CP element group try1_CP_1680_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(38) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_ZJ_357_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_ZJ_357_load_0_ack_1, ack => try1_CP_1680_elements(38)); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	33 
    -- CP-element group 39: successors 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	30 
    -- CP-element group 39: 	33 
    -- CP-element group 39: 	36 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_358_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_358_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_358_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_358_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_358_inst_ack_0, ack => try1_CP_1680_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_358_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_358_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_358_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(40) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_358_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_358_inst_ack_1, ack => try1_CP_1680_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	43 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/type_cast_363_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/type_cast_363_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/type_cast_363_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(41) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:type_cast_363_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(41), ack => type_cast_363_inst_req_0); -- 
    try1_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 24) := "try1_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(40) & try1_CP_1680_elements(43);
      gj_try1_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	51 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/type_cast_363_update_start_
      -- CP-element group 42: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/type_cast_363_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/type_cast_363_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(42) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:type_cast_363_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(42), ack => type_cast_363_inst_req_1); -- 
    try1_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(51);
      gj_try1_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	34 
    -- CP-element group 43: 	41 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/type_cast_363_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/type_cast_363_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/type_cast_363_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(43) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:type_cast_363_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_363_inst_ack_0, ack => try1_CP_1680_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/type_cast_363_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/type_cast_363_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/type_cast_363_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(44) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:type_cast_363_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_363_inst_ack_1, ack => try1_CP_1680_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: 	50 
    -- CP-element group 45: marked-predecessors 
    -- CP-element group 45: 	51 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	51 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/CONCAT_u1_u32_368_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/CONCAT_u1_u32_368_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/CONCAT_u1_u32_368_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(45) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:CONCAT_u1_u32_368_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(45), ack => CONCAT_u1_u32_368_inst_req_0); -- 
    try1_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 24) := "try1_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(44) & try1_CP_1680_elements(50) & try1_CP_1680_elements(51);
      gj_try1_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	55 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	52 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/CONCAT_u1_u32_368_update_start_
      -- CP-element group 46: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/CONCAT_u1_u32_368_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/CONCAT_u1_u32_368_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(46) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:CONCAT_u1_u32_368_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(46), ack => CONCAT_u1_u32_368_inst_req_1); -- 
    try1_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(55);
      gj_try1_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	9 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	49 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (5) 
      -- CP-element group 47: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_Sample/word_access_start/$entry
      -- CP-element group 47: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_Sample/word_access_start/word_0/$entry
      -- CP-element group 47: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(47) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_one_366_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(47), ack => LOAD_one_366_load_0_req_0); -- 
    try1_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 24) := "try1_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(9) & try1_CP_1680_elements(49);
      gj_try1_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: marked-predecessors 
    -- CP-element group 48: 	51 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (5) 
      -- CP-element group 48: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_update_start_
      -- CP-element group 48: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_Update/word_access_complete/$entry
      -- CP-element group 48: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_Update/word_access_complete/word_0/$entry
      -- CP-element group 48: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(48) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_one_366_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(48), ack => LOAD_one_366_load_0_req_1); -- 
    try1_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(51);
      gj_try1_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: marked-successors 
    -- CP-element group 49: 	47 
    -- CP-element group 49:  members (5) 
      -- CP-element group 49: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_Sample/word_access_start/$exit
      -- CP-element group 49: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_Sample/word_access_start/word_0/$exit
      -- CP-element group 49: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(49) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_one_366_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_one_366_load_0_ack_0, ack => try1_CP_1680_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	45 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_Update/word_access_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_Update/word_access_complete/word_0/$exit
      -- CP-element group 50: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_Update/word_access_complete/word_0/ca
      -- CP-element group 50: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_Update/LOAD_one_366_Merge/$entry
      -- CP-element group 50: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_Update/LOAD_one_366_Merge/$exit
      -- CP-element group 50: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_Update/LOAD_one_366_Merge/merge_req
      -- CP-element group 50: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/LOAD_one_366_Update/LOAD_one_366_Merge/merge_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(50) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_one_366_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_one_366_load_0_ack_1, ack => try1_CP_1680_elements(50)); -- 
    -- CP-element group 51:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	45 
    -- CP-element group 51: successors 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	42 
    -- CP-element group 51: 	45 
    -- CP-element group 51: 	48 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/CONCAT_u1_u32_368_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/CONCAT_u1_u32_368_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/CONCAT_u1_u32_368_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(51) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:CONCAT_u1_u32_368_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u1_u32_368_inst_ack_0, ack => try1_CP_1680_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	46 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/CONCAT_u1_u32_368_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/CONCAT_u1_u32_368_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/CONCAT_u1_u32_368_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(52) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:CONCAT_u1_u32_368_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u1_u32_368_inst_ack_1, ack => try1_CP_1680_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	55 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/call_stmt_373_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/call_stmt_373_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/call_stmt_373_Sample/crr
      -- 
    -- logger for CP element group try1_CP_1680_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(53) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:call_stmt_373_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(53), ack => call_stmt_373_call_req_0); -- 
    try1_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 24) := "try1_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(52) & try1_CP_1680_elements(55);
      gj_try1_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	87 
    -- CP-element group 54: 	91 
    -- CP-element group 54: 	59 
    -- CP-element group 54: 	63 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/call_stmt_373_update_start_
      -- CP-element group 54: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/call_stmt_373_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/call_stmt_373_Update/ccr
      -- 
    -- logger for CP element group try1_CP_1680_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(54) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:call_stmt_373_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_1888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(54), ack => call_stmt_373_call_req_1); -- 
    try1_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= try1_CP_1680_elements(87) & try1_CP_1680_elements(91) & try1_CP_1680_elements(59) & try1_CP_1680_elements(63);
      gj_try1_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: marked-successors 
    -- CP-element group 55: 	46 
    -- CP-element group 55: 	53 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/call_stmt_373_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/call_stmt_373_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/call_stmt_373_Sample/cra
      -- 
    -- logger for CP element group try1_CP_1680_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(55) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:call_stmt_373_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_373_call_ack_0, ack => try1_CP_1680_elements(55)); -- 
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	85 
    -- CP-element group 56: 	89 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	61 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/call_stmt_373_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/call_stmt_373_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/call_stmt_373_Update/cca
      -- 
    -- logger for CP element group try1_CP_1680_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(56) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:call_stmt_373_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_373_call_ack_1, ack => try1_CP_1680_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	59 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_376_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_376_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_376_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(57) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_376_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(57), ack => slice_376_inst_req_0); -- 
    try1_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 24) := "try1_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(56) & try1_CP_1680_elements(59);
      gj_try1_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	83 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_376_update_start_
      -- CP-element group 58: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_376_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_376_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(58) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_376_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(58), ack => slice_376_inst_req_1); -- 
    try1_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(83);
      gj_try1_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	54 
    -- CP-element group 59: 	57 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_376_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_376_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_376_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(59) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_376_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_376_inst_ack_0, ack => try1_CP_1680_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	81 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_376_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_376_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_376_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(60) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_376_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_376_inst_ack_1, ack => try1_CP_1680_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	56 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_380_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_380_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_380_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(61) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_380_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(61), ack => slice_380_inst_req_0); -- 
    try1_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 24) := "try1_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(56) & try1_CP_1680_elements(63);
      gj_try1_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	75 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_380_update_start_
      -- CP-element group 62: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_380_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_380_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(62) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_380_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(62), ack => slice_380_inst_req_1); -- 
    try1_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(75);
      gj_try1_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	54 
    -- CP-element group 63: 	61 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_380_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_380_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_380_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(63) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_380_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_380_inst_ack_0, ack => try1_CP_1680_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	73 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_380_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_380_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_380_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(64) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_380_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_380_inst_ack_1, ack => try1_CP_1680_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	15 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_385_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_385_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_385_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(65) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_385_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(65), ack => ADD_u12_u12_385_inst_req_0); -- 
    try1_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 24) := "try1_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(15) & try1_CP_1680_elements(67);
      gj_try1_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	79 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_385_update_start_
      -- CP-element group 66: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_385_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_385_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(66) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_385_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(66), ack => ADD_u12_u12_385_inst_req_1); -- 
    try1_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(79);
      gj_try1_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	13 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_385_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_385_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_385_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(67) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_385_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_385_inst_ack_0, ack => try1_CP_1680_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	77 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_385_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_385_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_385_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(68) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_385_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_385_inst_ack_1, ack => try1_CP_1680_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	15 
    -- CP-element group 69: marked-predecessors 
    -- CP-element group 69: 	71 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_389_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_389_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_389_Sample/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(69) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_T_341_delayed_12_0_387_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(69), ack => W_T_341_delayed_12_0_387_inst_req_0); -- 
    try1_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 24) := "try1_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(15) & try1_CP_1680_elements(71);
      gj_try1_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	75 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_389_update_start_
      -- CP-element group 70: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_389_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_389_Update/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(70)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(70)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(70) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_T_341_delayed_12_0_387_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(70), ack => W_T_341_delayed_12_0_387_inst_req_1); -- 
    try1_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(75);
      gj_try1_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	13 
    -- CP-element group 71: 	69 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_389_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_389_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_389_Sample/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(71)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(71)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(71) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_T_341_delayed_12_0_387_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_T_341_delayed_12_0_387_inst_ack_0, ack => try1_CP_1680_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (29) 
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_389_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_389_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_389_Update/ack
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_word_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_root_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_offset_calculated
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_index_resized_0
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_index_scaled_0
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_index_computed_0
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_index_resize_0/$entry
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_index_resize_0/$exit
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_index_resize_0/index_resize_req
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_index_resize_0/index_resize_ack
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_index_scale_0/$entry
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_index_scale_0/$exit
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_index_scale_0/scale_rename_req
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_index_scale_0/scale_rename_ack
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_final_index_sum_regn/$entry
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_final_index_sum_regn/$exit
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_final_index_sum_regn/req
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_final_index_sum_regn/ack
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_base_plus_offset/$entry
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_base_plus_offset/$exit
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_base_plus_offset/sum_rename_req
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_base_plus_offset/sum_rename_ack
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_word_addrgen/$entry
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_word_addrgen/$exit
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_word_addrgen/root_register_req
      -- CP-element group 72: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(72)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(72)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(72) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_T_341_delayed_12_0_387_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_T_341_delayed_12_0_387_inst_ack_1, ack => try1_CP_1680_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	64 
    -- CP-element group 73: 	72 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	115 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (9) 
      -- CP-element group 73: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_Sample/array_obj_ref_391_Split/$entry
      -- CP-element group 73: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_Sample/array_obj_ref_391_Split/$exit
      -- CP-element group 73: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_Sample/array_obj_ref_391_Split/split_req
      -- CP-element group 73: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_Sample/array_obj_ref_391_Split/split_ack
      -- CP-element group 73: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(73)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(73)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(73) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_391_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(73), ack => array_obj_ref_391_store_0_req_0); -- 
    try1_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 24) := "try1_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(64) & try1_CP_1680_elements(72) & try1_CP_1680_elements(115);
      gj_try1_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_update_start_
      -- CP-element group 74: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_Update/word_access_complete/$entry
      -- CP-element group 74: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_Update/word_access_complete/word_0/$entry
      -- CP-element group 74: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(74)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(74)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(74) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_391_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(74), ack => array_obj_ref_391_store_0_req_1); -- 
    try1_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(76);
      gj_try1_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	122 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	62 
    -- CP-element group 75: 	70 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_Sample/word_access_start/$exit
      -- CP-element group 75: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_Sample/word_access_start/word_0/$exit
      -- CP-element group 75: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(75)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(75)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(75) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_391_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_391_store_0_ack_0, ack => try1_CP_1680_elements(75)); -- 
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	125 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	74 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_Update/word_access_complete/$exit
      -- CP-element group 76: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_Update/word_access_complete/word_0/$exit
      -- CP-element group 76: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(76)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(76)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(76) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_391_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_391_store_0_ack_1, ack => try1_CP_1680_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	68 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	79 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_396_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_396_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_396_Sample/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(77)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(77)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(77) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_TT_345_delayed_11_0_394_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_2015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(77), ack => W_TT_345_delayed_11_0_394_inst_req_0); -- 
    try1_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 24) := "try1_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(68) & try1_CP_1680_elements(79);
      gj_try1_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	83 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_396_update_start_
      -- CP-element group 78: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_396_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_396_Update/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(78)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(78)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(78) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_TT_345_delayed_11_0_394_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_2020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(78), ack => W_TT_345_delayed_11_0_394_inst_req_1); -- 
    try1_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(83);
      gj_try1_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: 	66 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_396_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_396_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_396_Sample/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(79)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(79)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(79) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_TT_345_delayed_11_0_394_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_TT_345_delayed_11_0_394_inst_ack_0, ack => try1_CP_1680_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (29) 
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_396_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_396_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_396_Update/ack
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_word_address_calculated
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_root_address_calculated
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_offset_calculated
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_index_resized_0
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_index_scaled_0
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_index_computed_0
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_index_resize_0/$entry
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_index_resize_0/$exit
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_index_resize_0/index_resize_req
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_index_resize_0/index_resize_ack
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_index_scale_0/$entry
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_index_scale_0/$exit
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_index_scale_0/scale_rename_req
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_index_scale_0/scale_rename_ack
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_final_index_sum_regn/$entry
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_final_index_sum_regn/$exit
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_final_index_sum_regn/req
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_final_index_sum_regn/ack
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_base_plus_offset/$entry
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_base_plus_offset/$exit
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_base_plus_offset/sum_rename_req
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_base_plus_offset/sum_rename_ack
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_word_addrgen/$entry
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_word_addrgen/$exit
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_word_addrgen/root_register_req
      -- CP-element group 80: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(80)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(80)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(80) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_TT_345_delayed_11_0_394_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_TT_345_delayed_11_0_394_inst_ack_1, ack => try1_CP_1680_elements(80)); -- 
    -- CP-element group 81:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	122 
    -- CP-element group 81: 	80 
    -- CP-element group 81: 	60 
    -- CP-element group 81: marked-predecessors 
    -- CP-element group 81: 	83 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (9) 
      -- CP-element group 81: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_Sample/array_obj_ref_398_Split/$entry
      -- CP-element group 81: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_Sample/array_obj_ref_398_Split/$exit
      -- CP-element group 81: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_Sample/array_obj_ref_398_Split/split_req
      -- CP-element group 81: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_Sample/array_obj_ref_398_Split/split_ack
      -- CP-element group 81: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_Sample/word_access_start/$entry
      -- CP-element group 81: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_Sample/word_access_start/word_0/$entry
      -- CP-element group 81: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(81)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(81)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(81) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_398_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(81), ack => array_obj_ref_398_store_0_req_0); -- 
    try1_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 24) := "try1_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= try1_CP_1680_elements(122) & try1_CP_1680_elements(80) & try1_CP_1680_elements(60) & try1_CP_1680_elements(83);
      gj_try1_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: marked-predecessors 
    -- CP-element group 82: 	84 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (5) 
      -- CP-element group 82: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_update_start_
      -- CP-element group 82: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_Update/word_access_complete/$entry
      -- CP-element group 82: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_Update/word_access_complete/word_0/$entry
      -- CP-element group 82: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(82)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(82)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(82) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_398_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(82), ack => array_obj_ref_398_store_0_req_1); -- 
    try1_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(84);
      gj_try1_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	123 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	78 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	58 
    -- CP-element group 83:  members (5) 
      -- CP-element group 83: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_Sample/word_access_start/$exit
      -- CP-element group 83: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_Sample/word_access_start/word_0/$exit
      -- CP-element group 83: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(83)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(83)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(83) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_398_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_398_store_0_ack_0, ack => try1_CP_1680_elements(83)); -- 
    -- CP-element group 84:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	125 
    -- CP-element group 84: marked-successors 
    -- CP-element group 84: 	82 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_Update/word_access_complete/$exit
      -- CP-element group 84: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_Update/word_access_complete/word_0/$exit
      -- CP-element group 84: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(84)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(84)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(84) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_398_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_398_store_0_ack_1, ack => try1_CP_1680_elements(84)); -- 
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	56 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_403_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_403_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_403_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(85)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(85)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(85) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_403_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(85), ack => slice_403_inst_req_0); -- 
    try1_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 24) := "try1_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(56) & try1_CP_1680_elements(87);
      gj_try1_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: marked-predecessors 
    -- CP-element group 86: 	115 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_403_update_start_
      -- CP-element group 86: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_403_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_403_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(86)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(86)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(86) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_403_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(86), ack => slice_403_inst_req_1); -- 
    try1_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(115);
      gj_try1_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	54 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_403_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_403_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_403_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(87)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(87)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(87) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_403_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_403_inst_ack_0, ack => try1_CP_1680_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	113 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_403_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_403_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_403_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(88)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(88)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(88) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_403_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_403_inst_ack_1, ack => try1_CP_1680_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	56 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_407_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_407_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_407_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(89)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(89)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(89) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_407_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(89), ack => slice_407_inst_req_0); -- 
    try1_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 24) := "try1_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(56) & try1_CP_1680_elements(91);
      gj_try1_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	107 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_407_update_start_
      -- CP-element group 90: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_407_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_407_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(90)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(90)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(90) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_407_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(90), ack => slice_407_inst_req_1); -- 
    try1_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(107);
      gj_try1_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	54 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_407_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_407_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_407_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(91)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(91)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(91) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_407_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_407_inst_ack_0, ack => try1_CP_1680_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	105 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_407_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_407_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/slice_407_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(92)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(92)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(92) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_407_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_407_inst_ack_1, ack => try1_CP_1680_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	15 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	95 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_412_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_412_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_412_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(93)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(93)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(93) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_412_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(93), ack => ADD_u12_u12_412_inst_req_0); -- 
    try1_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 24) := "try1_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(15) & try1_CP_1680_elements(95);
      gj_try1_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	103 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_412_update_start_
      -- CP-element group 94: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_412_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_412_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(94)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(94)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(94) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_412_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(94), ack => ADD_u12_u12_412_inst_req_1); -- 
    try1_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(103);
      gj_try1_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	13 
    -- CP-element group 95: 	93 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_412_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_412_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_412_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(95)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(95)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(95) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_412_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_412_inst_ack_0, ack => try1_CP_1680_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	101 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_412_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_412_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_412_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(96)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(96)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(96) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_412_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_412_inst_ack_1, ack => try1_CP_1680_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	15 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	99 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_417_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_417_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_417_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(97)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(97)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(97) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_417_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(97), ack => ADD_u12_u12_417_inst_req_0); -- 
    try1_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 24) := "try1_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(15) & try1_CP_1680_elements(99);
      gj_try1_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	111 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_417_update_start_
      -- CP-element group 98: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_417_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_417_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(98)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(98)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(98) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_417_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(98), ack => ADD_u12_u12_417_inst_req_1); -- 
    try1_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(111);
      gj_try1_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	13 
    -- CP-element group 99: 	97 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_417_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_417_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_417_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(99)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(99)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(99) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_417_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_417_inst_ack_0, ack => try1_CP_1680_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	109 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_417_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_417_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_417_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(100)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(100)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(100) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_417_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_417_inst_ack_1, ack => try1_CP_1680_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	96 
    -- CP-element group 101: marked-predecessors 
    -- CP-element group 101: 	103 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_421_sample_start_
      -- CP-element group 101: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_421_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_421_Sample/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(101)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(101)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(101) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_TTT_367_delayed_11_0_419_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_2147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(101), ack => W_TTT_367_delayed_11_0_419_inst_req_0); -- 
    try1_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(96) & try1_CP_1680_elements(103);
      gj_try1_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: marked-predecessors 
    -- CP-element group 102: 	107 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_421_update_start_
      -- CP-element group 102: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_421_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_421_Update/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(102)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(102)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(102) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_TTT_367_delayed_11_0_419_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_2152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(102), ack => W_TTT_367_delayed_11_0_419_inst_req_1); -- 
    try1_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(107);
      gj_try1_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: marked-successors 
    -- CP-element group 103: 	94 
    -- CP-element group 103: 	101 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_421_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_421_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_421_Sample/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(103)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(103)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(103) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_TTT_367_delayed_11_0_419_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_TTT_367_delayed_11_0_419_inst_ack_0, ack => try1_CP_1680_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (29) 
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_421_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_421_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_421_Update/ack
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_word_address_calculated
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_root_address_calculated
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_offset_calculated
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_index_resized_0
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_index_scaled_0
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_index_computed_0
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_index_resize_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_index_resize_0/$exit
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_index_resize_0/index_resize_req
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_index_resize_0/index_resize_ack
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_index_scale_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_index_scale_0/$exit
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_index_scale_0/scale_rename_req
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_index_scale_0/scale_rename_ack
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_final_index_sum_regn/$entry
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_final_index_sum_regn/$exit
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_final_index_sum_regn/req
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_final_index_sum_regn/ack
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_base_plus_offset/$entry
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_base_plus_offset/$exit
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_base_plus_offset/sum_rename_req
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_base_plus_offset/sum_rename_ack
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_word_addrgen/$entry
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_word_addrgen/$exit
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_word_addrgen/root_register_req
      -- CP-element group 104: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(104)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(104)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(104) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_TTT_367_delayed_11_0_419_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_TTT_367_delayed_11_0_419_inst_ack_1, ack => try1_CP_1680_elements(104)); -- 
    -- CP-element group 105:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	123 
    -- CP-element group 105: 	92 
    -- CP-element group 105: 	104 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	107 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (9) 
      -- CP-element group 105: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_Sample/array_obj_ref_423_Split/$entry
      -- CP-element group 105: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_Sample/array_obj_ref_423_Split/$exit
      -- CP-element group 105: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_Sample/array_obj_ref_423_Split/split_req
      -- CP-element group 105: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_Sample/array_obj_ref_423_Split/split_ack
      -- CP-element group 105: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_Sample/word_access_start/$entry
      -- CP-element group 105: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_Sample/word_access_start/word_0/$entry
      -- CP-element group 105: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(105)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(105)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(105) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_423_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(105), ack => array_obj_ref_423_store_0_req_0); -- 
    try1_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= try1_CP_1680_elements(123) & try1_CP_1680_elements(92) & try1_CP_1680_elements(104) & try1_CP_1680_elements(107);
      gj_try1_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: marked-predecessors 
    -- CP-element group 106: 	108 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (5) 
      -- CP-element group 106: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_update_start_
      -- CP-element group 106: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_Update/word_access_complete/$entry
      -- CP-element group 106: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_Update/word_access_complete/word_0/$entry
      -- CP-element group 106: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(106)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(106)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(106) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_423_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(106), ack => array_obj_ref_423_store_0_req_1); -- 
    try1_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(108);
      gj_try1_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	124 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	102 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	90 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_Sample/word_access_start/$exit
      -- CP-element group 107: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_Sample/word_access_start/word_0/$exit
      -- CP-element group 107: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(107)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(107)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(107) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_423_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_423_store_0_ack_0, ack => try1_CP_1680_elements(107)); -- 
    -- CP-element group 108:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	125 
    -- CP-element group 108: marked-successors 
    -- CP-element group 108: 	106 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_Update/word_access_complete/$exit
      -- CP-element group 108: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_Update/word_access_complete/word_0/$exit
      -- CP-element group 108: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(108)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(108)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(108) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_423_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_423_store_0_ack_1, ack => try1_CP_1680_elements(108)); -- 
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	100 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	111 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_428_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_428_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_428_Sample/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(109)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(109)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(109) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_TTTT_371_delayed_11_0_426_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_2223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(109), ack => W_TTTT_371_delayed_11_0_426_inst_req_0); -- 
    try1_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(100) & try1_CP_1680_elements(111);
      gj_try1_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	115 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_428_update_start_
      -- CP-element group 110: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_428_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_428_Update/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(110)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(110)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(110) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_TTTT_371_delayed_11_0_426_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_2228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(110), ack => W_TTTT_371_delayed_11_0_426_inst_req_1); -- 
    try1_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(115);
      gj_try1_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: marked-successors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	98 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_428_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_428_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_428_Sample/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(111)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(111)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(111) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_TTTT_371_delayed_11_0_426_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_TTTT_371_delayed_11_0_426_inst_ack_0, ack => try1_CP_1680_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (29) 
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_base_plus_offset/sum_rename_ack
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_word_addrgen/root_register_ack
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_word_addrgen/$entry
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_base_plus_offset/$entry
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_base_plus_offset/$exit
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_word_addrgen/$exit
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_base_plus_offset/sum_rename_req
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_word_addrgen/root_register_req
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_428_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_428_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/assign_stmt_428_Update/ack
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_word_address_calculated
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_root_address_calculated
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_offset_calculated
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_index_resized_0
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_index_scaled_0
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_index_computed_0
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_index_resize_0/$entry
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_index_resize_0/$exit
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_index_resize_0/index_resize_req
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_index_resize_0/index_resize_ack
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_index_scale_0/$entry
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_index_scale_0/$exit
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_index_scale_0/scale_rename_req
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_index_scale_0/scale_rename_ack
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_final_index_sum_regn/$entry
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_final_index_sum_regn/$exit
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_final_index_sum_regn/req
      -- CP-element group 112: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_final_index_sum_regn/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(112)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(112)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(112) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_TTTT_371_delayed_11_0_426_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_TTTT_371_delayed_11_0_426_inst_ack_1, ack => try1_CP_1680_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: 	124 
    -- CP-element group 113: 	88 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	115 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (9) 
      -- CP-element group 113: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_Sample/word_access_start/$entry
      -- CP-element group 113: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_Sample/word_access_start/word_0/rr
      -- CP-element group 113: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_Sample/array_obj_ref_430_Split/$exit
      -- CP-element group 113: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_Sample/word_access_start/word_0/$entry
      -- CP-element group 113: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_Sample/array_obj_ref_430_Split/split_req
      -- CP-element group 113: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_Sample/array_obj_ref_430_Split/split_ack
      -- CP-element group 113: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_Sample/array_obj_ref_430_Split/$entry
      -- CP-element group 113: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_sample_start_
      -- 
    -- logger for CP element group try1_CP_1680_elements(113)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(113)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(113) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_430_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(113), ack => array_obj_ref_430_store_0_req_0); -- 
    try1_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= try1_CP_1680_elements(112) & try1_CP_1680_elements(124) & try1_CP_1680_elements(88) & try1_CP_1680_elements(115);
      gj_try1_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	116 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (5) 
      -- CP-element group 114: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_Update/word_access_complete/$entry
      -- CP-element group 114: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_Update/word_access_complete/word_0/$entry
      -- CP-element group 114: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_Update/word_access_complete/word_0/cr
      -- CP-element group 114: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_update_start_
      -- 
    -- logger for CP element group try1_CP_1680_elements(114)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(114)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(114) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_430_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(114), ack => array_obj_ref_430_store_0_req_1); -- 
    try1_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(116);
      gj_try1_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	125 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	110 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	86 
    -- CP-element group 115: 	73 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_Sample/word_access_start/word_0/ra
      -- CP-element group 115: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_Sample/word_access_start/$exit
      -- CP-element group 115: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_Sample/word_access_start/word_0/$exit
      -- CP-element group 115: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ring_reenable_memory_space_4
      -- 
    -- logger for CP element group try1_CP_1680_elements(115)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(115)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(115) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_430_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_430_store_0_ack_0, ack => try1_CP_1680_elements(115)); -- 
    -- CP-element group 116:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	125 
    -- CP-element group 116: marked-successors 
    -- CP-element group 116: 	114 
    -- CP-element group 116:  members (5) 
      -- CP-element group 116: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_Update/word_access_complete/$exit
      -- CP-element group 116: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_Update/word_access_complete/word_0/ca
      -- CP-element group 116: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_Update/word_access_complete/word_0/$exit
      -- CP-element group 116: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_430_update_completed_
      -- 
    -- logger for CP element group try1_CP_1680_elements(116)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(116)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(116) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_430_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_430_store_0_ack_1, ack => try1_CP_1680_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	15 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	119 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_436_sample_start_
      -- CP-element group 117: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_436_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_436_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(117)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(117)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(117) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_436_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(117), ack => ADD_u12_u12_436_inst_req_0); -- 
    try1_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(15) & try1_CP_1680_elements(119);
      gj_try1_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	14 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	120 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_436_update_start_
      -- CP-element group 118: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_436_Update/$entry
      -- CP-element group 118: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_436_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(118)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(118)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(118) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_436_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(118), ack => ADD_u12_u12_436_inst_req_1); -- 
    try1_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(14) & try1_CP_1680_elements(120);
      gj_try1_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: successors 
    -- CP-element group 119: marked-successors 
    -- CP-element group 119: 	13 
    -- CP-element group 119: 	117 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_436_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_436_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_436_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(119)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(119)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(119) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_436_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_436_inst_ack_0, ack => try1_CP_1680_elements(119)); -- 
    -- CP-element group 120:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	10 
    -- CP-element group 120: marked-successors 
    -- CP-element group 120: 	12 
    -- CP-element group 120: 	118 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_436_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_436_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/ADD_u12_u12_436_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(120)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(120)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(120) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_436_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_436_inst_ack_1, ack => try1_CP_1680_elements(120)); -- 
    -- CP-element group 121:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	9 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	10 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group try1_CP_1680_elements(121)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(121)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(121) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(121) is a control-delay.
    cp_element_121_delay: control_delay_element  generic map(name => " 121_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(9), ack => try1_CP_1680_elements(121), clk => clk, reset =>reset);
    -- CP-element group 122:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	75 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	81 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_391_array_obj_ref_398_delay
      -- 
    -- logger for CP element group try1_CP_1680_elements(122)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(122)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(122) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(122) is a control-delay.
    cp_element_122_delay: control_delay_element  generic map(name => " 122_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(75), ack => try1_CP_1680_elements(122), clk => clk, reset =>reset);
    -- CP-element group 123:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	83 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	105 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_398_array_obj_ref_423_delay
      -- 
    -- logger for CP element group try1_CP_1680_elements(123)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(123)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(123) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(123) is a control-delay.
    cp_element_123_delay: control_delay_element  generic map(name => " 123_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(83), ack => try1_CP_1680_elements(123), clk => clk, reset =>reset);
    -- CP-element group 124:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	107 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	113 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/array_obj_ref_423_array_obj_ref_430_delay
      -- 
    -- logger for CP element group try1_CP_1680_elements(124)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(124)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(124) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(124) is a control-delay.
    cp_element_124_delay: control_delay_element  generic map(name => " 124_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(107), ack => try1_CP_1680_elements(124), clk => clk, reset =>reset);
    -- CP-element group 125:  join  transition  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	76 
    -- CP-element group 125: 	108 
    -- CP-element group 125: 	115 
    -- CP-element group 125: 	116 
    -- CP-element group 125: 	84 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	6 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_343/do_while_stmt_344/do_while_stmt_344_loop_body/$exit
      -- 
    -- logger for CP element group try1_CP_1680_elements(125)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(125)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(125) fired."); 
        -- 
      end if; --
    end process; 
    try1_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= try1_CP_1680_elements(76) & try1_CP_1680_elements(108) & try1_CP_1680_elements(115) & try1_CP_1680_elements(116) & try1_CP_1680_elements(84);
      gj_try1_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	5 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_343/do_while_stmt_344/loop_exit/$exit
      -- CP-element group 126: 	 branch_block_stmt_343/do_while_stmt_344/loop_exit/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(126)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(126)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(126) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:do_while_stmt_344_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_344_branch_ack_0, ack => try1_CP_1680_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	5 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_343/do_while_stmt_344/loop_taken/$exit
      -- CP-element group 127: 	 branch_block_stmt_343/do_while_stmt_344/loop_taken/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(127)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(127)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(127) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:do_while_stmt_344_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_344_branch_ack_1, ack => try1_CP_1680_elements(127)); -- 
    -- CP-element group 128:  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	3 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	1 
    -- CP-element group 128:  members (1) 
      -- CP-element group 128: 	 branch_block_stmt_343/do_while_stmt_344/$exit
      -- 
    -- logger for CP element group try1_CP_1680_elements(128)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(128)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(128) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(128) <= try1_CP_1680_elements(3);
    -- CP-element group 129:  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	527 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (5) 
      -- CP-element group 129: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_Sample/word_access_start/$exit
      -- CP-element group 129: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_Sample/word_access_start/word_0/$exit
      -- CP-element group 129: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(129)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(129)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(129) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:STORE_PJ_451_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_PJ_451_store_0_ack_0, ack => try1_CP_1680_elements(129)); -- 
    -- CP-element group 130:  transition  place  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	527 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (11) 
      -- CP-element group 130: 	 branch_block_stmt_443/branch_block_stmt_454__entry__
      -- CP-element group 130: 	 branch_block_stmt_443/assign_stmt_453__exit__
      -- CP-element group 130: 	 branch_block_stmt_443/branch_block_stmt_454/branch_block_stmt_454__entry__
      -- CP-element group 130: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455__entry__
      -- CP-element group 130: 	 branch_block_stmt_443/assign_stmt_453/$exit
      -- CP-element group 130: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_Update/word_access_complete/$exit
      -- CP-element group 130: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_Update/word_access_complete/word_0/$exit
      -- CP-element group 130: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_Update/word_access_complete/word_0/ca
      -- CP-element group 130: 	 branch_block_stmt_443/branch_block_stmt_454/$entry
      -- 
    -- logger for CP element group try1_CP_1680_elements(130)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(130)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(130) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:STORE_PJ_451_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_PJ_451_store_0_ack_1, ack => try1_CP_1680_elements(130)); -- 
    -- CP-element group 131:  branch  transition  place  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	291 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	512 
    -- CP-element group 131:  members (12) 
      -- CP-element group 131: 	 branch_block_stmt_443/branch_block_stmt_565__entry__
      -- CP-element group 131: 	 branch_block_stmt_443/branch_block_stmt_565/merge_stmt_566__entry__
      -- CP-element group 131: 	 branch_block_stmt_443/branch_block_stmt_454__exit__
      -- CP-element group 131: 	 branch_block_stmt_443/branch_block_stmt_454/branch_block_stmt_454__exit__
      -- CP-element group 131: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455__exit__
      -- CP-element group 131: 	 branch_block_stmt_443/branch_block_stmt_454/$exit
      -- CP-element group 131: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_565__entry__
      -- CP-element group 131: 	 branch_block_stmt_443/branch_block_stmt_565/$entry
      -- CP-element group 131: 	 branch_block_stmt_443/branch_block_stmt_565/merge_stmt_566_dead_link/$entry
      -- CP-element group 131: 	 branch_block_stmt_443/branch_block_stmt_565/merge_stmt_566__entry___PhiReq/$entry
      -- CP-element group 131: 	 branch_block_stmt_443/branch_block_stmt_565/merge_stmt_566__entry___PhiReq/phi_stmt_567/$entry
      -- CP-element group 131: 	 branch_block_stmt_443/branch_block_stmt_565/merge_stmt_566__entry___PhiReq/phi_stmt_567/phi_stmt_567_sources/$entry
      -- 
    -- logger for CP element group try1_CP_1680_elements(131)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(131)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(131) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(131) <= try1_CP_1680_elements(291);
    -- CP-element group 132:  transition  place  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	138 
    -- CP-element group 132:  members (2) 
      -- CP-element group 132: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455__entry__
      -- CP-element group 132: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/$entry
      -- 
    -- logger for CP element group try1_CP_1680_elements(132)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(132)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(132) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(132) <= try1_CP_1680_elements(130);
    -- CP-element group 133:  merge  place  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	291 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455__exit__
      -- 
    -- logger for CP element group try1_CP_1680_elements(133)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(133)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(133) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(133) is bound as output of CP function.
    -- CP-element group 134:  merge  place  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (1) 
      -- CP-element group 134: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/loop_back
      -- 
    -- logger for CP element group try1_CP_1680_elements(134)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(134)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(134) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(134) is bound as output of CP function.
    -- CP-element group 135:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	140 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	289 
    -- CP-element group 135: 	290 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/condition_done
      -- CP-element group 135: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/loop_exit/$entry
      -- CP-element group 135: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/loop_taken/$entry
      -- 
    -- logger for CP element group try1_CP_1680_elements(135)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(135)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(135) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(135) <= try1_CP_1680_elements(140);
    -- CP-element group 136:  branch  place  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	288 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/loop_body_done
      -- 
    -- logger for CP element group try1_CP_1680_elements(136)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(136)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(136) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(136) <= try1_CP_1680_elements(288);
    -- CP-element group 137:  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	146 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group try1_CP_1680_elements(137)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(137)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(137) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(137) <= try1_CP_1680_elements(134);
    -- CP-element group 138:  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	132 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	148 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group try1_CP_1680_elements(138)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(138)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(138) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(138) <= try1_CP_1680_elements(132);
    -- CP-element group 139:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	163 
    -- CP-element group 139: 	142 
    -- CP-element group 139: 	143 
    -- CP-element group 139: 	201 
    -- CP-element group 139: 	269 
    -- CP-element group 139: 	275 
    -- CP-element group 139: 	279 
    -- CP-element group 139: 	207 
    -- CP-element group 139: 	173 
    -- CP-element group 139: 	233 
    -- CP-element group 139: 	241 
    -- CP-element group 139:  members (16) 
      -- CP-element group 139: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_root_address_calculated
      -- CP-element group 139: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_word_address_calculated
      -- CP-element group 139: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_root_address_calculated
      -- CP-element group 139: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_word_address_calculated
      -- CP-element group 139: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/$entry
      -- CP-element group 139: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/loop_body_start
      -- CP-element group 139: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_word_address_calculated
      -- CP-element group 139: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_root_address_calculated
      -- CP-element group 139: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_word_address_calculated
      -- CP-element group 139: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_root_address_calculated
      -- CP-element group 139: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_word_address_calculated
      -- CP-element group 139: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_root_address_calculated
      -- CP-element group 139: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_word_address_calculated
      -- CP-element group 139: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_root_address_calculated
      -- CP-element group 139: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_word_address_calculated
      -- CP-element group 139: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_root_address_calculated
      -- 
    -- logger for CP element group try1_CP_1680_elements(139)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(139)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(139) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(139) is bound as output of CP function.
    -- CP-element group 140:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	145 
    -- CP-element group 140: 	266 
    -- CP-element group 140: 	279 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	135 
    -- CP-element group 140:  members (1) 
      -- CP-element group 140: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/condition_evaluated
      -- 
    -- logger for CP element group try1_CP_1680_elements(140)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(140)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(140) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:do_while_stmt_455_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_2394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(140), ack => do_while_stmt_455_branch_req_0); -- 
    try1_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(145) & try1_CP_1680_elements(266) & try1_CP_1680_elements(279);
      gj_try1_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	142 
    -- CP-element group 141: marked-predecessors 
    -- CP-element group 141: 	145 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (2) 
      -- CP-element group 141: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/aggregated_phi_sample_req
      -- CP-element group 141: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/phi_stmt_457_sample_start__ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(141)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(141)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(141) fired."); 
        -- 
      end if; --
    end process; 
    try1_cp_element_group_141: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_141"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(142) & try1_CP_1680_elements(145);
      gj_try1_cp_element_group_141 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 142:  join  transition  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	139 
    -- CP-element group 142: marked-predecessors 
    -- CP-element group 142: 	144 
    -- CP-element group 142: 	266 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	141 
    -- CP-element group 142:  members (1) 
      -- CP-element group 142: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/phi_stmt_457_sample_start_
      -- 
    -- logger for CP element group try1_CP_1680_elements(142)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(142)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(142) fired."); 
        -- 
      end if; --
    end process; 
    try1_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(139) & try1_CP_1680_elements(144) & try1_CP_1680_elements(266);
      gj_try1_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	139 
    -- CP-element group 143: marked-predecessors 
    -- CP-element group 143: 	161 
    -- CP-element group 143: 	145 
    -- CP-element group 143: 	265 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/aggregated_phi_update_req
      -- CP-element group 143: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/phi_stmt_457_update_start_
      -- CP-element group 143: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/phi_stmt_457_update_start__ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(143)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(143)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(143) fired."); 
        -- 
      end if; --
    end process; 
    try1_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= try1_CP_1680_elements(139) & try1_CP_1680_elements(161) & try1_CP_1680_elements(145) & try1_CP_1680_elements(265);
      gj_try1_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	264 
    -- CP-element group 144: marked-successors 
    -- CP-element group 144: 	142 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/aggregated_phi_sample_ack
      -- CP-element group 144: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/phi_stmt_457_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/phi_stmt_457_sample_completed__ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(144)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(144)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(144) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(144) is bound as output of CP function.
    -- CP-element group 145:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	159 
    -- CP-element group 145: 	140 
    -- CP-element group 145: 	263 
    -- CP-element group 145: marked-successors 
    -- CP-element group 145: 	141 
    -- CP-element group 145: 	143 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/aggregated_phi_update_ack
      -- CP-element group 145: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/phi_stmt_457_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/phi_stmt_457_update_completed__ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(145)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(145)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(145) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(145) is bound as output of CP function.
    -- CP-element group 146:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	137 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (1) 
      -- CP-element group 146: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/phi_stmt_457_loopback_trigger
      -- 
    -- logger for CP element group try1_CP_1680_elements(146)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(146)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(146) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(146) <= try1_CP_1680_elements(137);
    -- CP-element group 147:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/phi_stmt_457_loopback_sample_req
      -- CP-element group 147: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/phi_stmt_457_loopback_sample_req_ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(147)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(147)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(147) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:phi_stmt_457_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_457_loopback_sample_req_2409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_457_loopback_sample_req_2409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(147), ack => phi_stmt_457_req_1); -- 
    -- Element group try1_CP_1680_elements(147) is bound as output of CP function.
    -- CP-element group 148:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	138 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (1) 
      -- CP-element group 148: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/phi_stmt_457_entry_trigger
      -- 
    -- logger for CP element group try1_CP_1680_elements(148)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(148)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(148) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(148) <= try1_CP_1680_elements(138);
    -- CP-element group 149:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (2) 
      -- CP-element group 149: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/phi_stmt_457_entry_sample_req
      -- CP-element group 149: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/phi_stmt_457_entry_sample_req_ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(149)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(149)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(149) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:phi_stmt_457_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_457_entry_sample_req_2412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_457_entry_sample_req_2412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(149), ack => phi_stmt_457_req_0); -- 
    -- Element group try1_CP_1680_elements(149) is bound as output of CP function.
    -- CP-element group 150:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: successors 
    -- CP-element group 150:  members (2) 
      -- CP-element group 150: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/phi_stmt_457_phi_mux_ack
      -- CP-element group 150: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/phi_stmt_457_phi_mux_ack_ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(150)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(150)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(150) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:phi_stmt_457_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_457_phi_mux_ack_2415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_457_ack_0, ack => try1_CP_1680_elements(150)); -- 
    -- CP-element group 151:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (4) 
      -- CP-element group 151: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_460_sample_start__ps
      -- CP-element group 151: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_460_sample_completed__ps
      -- CP-element group 151: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_460_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_460_sample_completed_
      -- 
    -- logger for CP element group try1_CP_1680_elements(151)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(151)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(151) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(151) is bound as output of CP function.
    -- CP-element group 152:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (2) 
      -- CP-element group 152: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_460_update_start__ps
      -- CP-element group 152: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_460_update_start_
      -- 
    -- logger for CP element group try1_CP_1680_elements(152)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(152)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(152) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(152) is bound as output of CP function.
    -- CP-element group 153:  join  transition  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	154 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (1) 
      -- CP-element group 153: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_460_update_completed__ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(153)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(153)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(153) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(153) <= try1_CP_1680_elements(154);
    -- CP-element group 154:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	153 
    -- CP-element group 154:  members (1) 
      -- CP-element group 154: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_460_update_completed_
      -- 
    -- logger for CP element group try1_CP_1680_elements(154)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(154)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(154) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(154) is a control-delay.
    cp_element_154_delay: control_delay_element  generic map(name => " 154_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(152), ack => try1_CP_1680_elements(154), clk => clk, reset =>reset);
    -- CP-element group 155:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (4) 
      -- CP-element group 155: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/R_NJ_461_sample_start__ps
      -- CP-element group 155: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/R_NJ_461_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/R_NJ_461_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/R_NJ_461_Sample/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(155)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(155)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(155) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NJ_554_461_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_2436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(155), ack => NJ_554_461_buf_req_0); -- 
    -- Element group try1_CP_1680_elements(155) is bound as output of CP function.
    -- CP-element group 156:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (4) 
      -- CP-element group 156: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/R_NJ_461_update_start__ps
      -- CP-element group 156: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/R_NJ_461_update_start_
      -- CP-element group 156: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/R_NJ_461_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/R_NJ_461_Update/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(156)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(156)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(156) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NJ_554_461_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_2441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(156), ack => NJ_554_461_buf_req_1); -- 
    -- Element group try1_CP_1680_elements(156) is bound as output of CP function.
    -- CP-element group 157:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157:  members (4) 
      -- CP-element group 157: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/R_NJ_461_sample_completed__ps
      -- CP-element group 157: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/R_NJ_461_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/R_NJ_461_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/R_NJ_461_Sample/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(157)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(157)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(157) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NJ_554_461_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NJ_554_461_buf_ack_0, ack => try1_CP_1680_elements(157)); -- 
    -- CP-element group 158:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (4) 
      -- CP-element group 158: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/R_NJ_461_update_completed__ps
      -- CP-element group 158: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/R_NJ_461_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/R_NJ_461_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/R_NJ_461_Update/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(158)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(158)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(158) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NJ_554_461_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NJ_554_461_buf_ack_1, ack => try1_CP_1680_elements(158)); -- 
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	145 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	161 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_465_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_465_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_465_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(159)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(159)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(159) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:type_cast_465_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(159), ack => type_cast_465_inst_req_0); -- 
    try1_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(145) & try1_CP_1680_elements(161);
      gj_try1_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	169 
    -- CP-element group 160: 	162 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_465_update_start_
      -- CP-element group 160: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_465_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_465_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(160)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(160)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(160) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:type_cast_465_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(160), ack => type_cast_465_inst_req_1); -- 
    try1_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(169) & try1_CP_1680_elements(162);
      gj_try1_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: 	143 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_465_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_465_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_465_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(161)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(161)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(161) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:type_cast_465_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_465_inst_ack_0, ack => try1_CP_1680_elements(161)); -- 
    -- CP-element group 162:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	167 
    -- CP-element group 162: marked-successors 
    -- CP-element group 162: 	160 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_465_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_465_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_465_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(162)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(162)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(162) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:type_cast_465_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_465_inst_ack_1, ack => try1_CP_1680_elements(162)); -- 
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	139 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_469_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_469_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_469_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(163)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(163)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(163) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:type_cast_469_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(163), ack => type_cast_469_inst_req_0); -- 
    try1_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(139) & try1_CP_1680_elements(165);
      gj_try1_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	166 
    -- CP-element group 164: 	181 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_469_update_start_
      -- CP-element group 164: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_469_Update/$entry
      -- CP-element group 164: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_469_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(164)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(164)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(164) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:type_cast_469_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(164), ack => type_cast_469_inst_req_1); -- 
    try1_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(166) & try1_CP_1680_elements(181);
      gj_try1_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	163 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_469_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_469_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_469_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(165)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(165)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(165) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:type_cast_469_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_469_inst_ack_0, ack => try1_CP_1680_elements(165)); -- 
    -- CP-element group 166:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	179 
    -- CP-element group 166: marked-successors 
    -- CP-element group 166: 	164 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_469_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_469_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/type_cast_469_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(166)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(166)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(166) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:type_cast_469_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_469_inst_ack_1, ack => try1_CP_1680_elements(166)); -- 
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	162 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	169 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_473_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_473_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_473_Sample/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(167)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(167)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(167) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_NJJ_415_delayed_2_0_471_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_2479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(167), ack => W_NJJ_415_delayed_2_0_471_inst_req_0); -- 
    try1_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(162) & try1_CP_1680_elements(169);
      gj_try1_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	177 
    -- CP-element group 168: 	170 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_473_update_start_
      -- CP-element group 168: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_473_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_473_Update/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(168)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(168)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(168) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_NJJ_415_delayed_2_0_471_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_2484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(168), ack => W_NJJ_415_delayed_2_0_471_inst_req_1); -- 
    try1_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(177) & try1_CP_1680_elements(170);
      gj_try1_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: marked-successors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: 	160 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_473_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_473_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_473_Sample/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(169)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(169)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(169) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_NJJ_415_delayed_2_0_471_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_NJJ_415_delayed_2_0_471_inst_ack_0, ack => try1_CP_1680_elements(169)); -- 
    -- CP-element group 170:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	168 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_473_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_473_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_473_Update/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(170)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(170)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(170) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_NJJ_415_delayed_2_0_471_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_NJJ_415_delayed_2_0_471_inst_ack_1, ack => try1_CP_1680_elements(170)); -- 
    -- CP-element group 171:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	176 
    -- CP-element group 171: 	170 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	177 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	177 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/CONCAT_u1_u32_477_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/CONCAT_u1_u32_477_Sample/$entry
      -- CP-element group 171: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/CONCAT_u1_u32_477_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(171)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(171)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(171) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:CONCAT_u1_u32_477_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(171), ack => CONCAT_u1_u32_477_inst_req_0); -- 
    try1_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(176) & try1_CP_1680_elements(170) & try1_CP_1680_elements(177);
      gj_try1_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	185 
    -- CP-element group 172: 	178 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	178 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/CONCAT_u1_u32_477_update_start_
      -- CP-element group 172: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/CONCAT_u1_u32_477_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/CONCAT_u1_u32_477_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(172)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(172)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(172) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:CONCAT_u1_u32_477_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(172), ack => CONCAT_u1_u32_477_inst_req_1); -- 
    try1_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(185) & try1_CP_1680_elements(178);
      gj_try1_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	139 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (5) 
      -- CP-element group 173: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_sample_start_
      -- CP-element group 173: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_Sample/$entry
      -- CP-element group 173: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_Sample/word_access_start/$entry
      -- CP-element group 173: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_Sample/word_access_start/word_0/$entry
      -- CP-element group 173: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(173)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(173)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(173) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_one_475_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(173), ack => LOAD_one_475_load_0_req_0); -- 
    try1_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(139) & try1_CP_1680_elements(175);
      gj_try1_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: marked-predecessors 
    -- CP-element group 174: 	176 
    -- CP-element group 174: 	177 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (5) 
      -- CP-element group 174: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_update_start_
      -- CP-element group 174: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_Update/$entry
      -- CP-element group 174: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_Update/word_access_complete/$entry
      -- CP-element group 174: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_Update/word_access_complete/word_0/$entry
      -- CP-element group 174: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(174)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(174)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(174) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_one_475_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(174), ack => LOAD_one_475_load_0_req_1); -- 
    try1_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(176) & try1_CP_1680_elements(177);
      gj_try1_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	173 
    -- CP-element group 175:  members (5) 
      -- CP-element group 175: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_Sample/word_access_start/$exit
      -- CP-element group 175: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_Sample/word_access_start/word_0/$exit
      -- CP-element group 175: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(175)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(175)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(175) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_one_475_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_one_475_load_0_ack_0, ack => try1_CP_1680_elements(175)); -- 
    -- CP-element group 176:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	171 
    -- CP-element group 176: marked-successors 
    -- CP-element group 176: 	174 
    -- CP-element group 176:  members (9) 
      -- CP-element group 176: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_Update/word_access_complete/$exit
      -- CP-element group 176: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_Update/word_access_complete/word_0/$exit
      -- CP-element group 176: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_Update/word_access_complete/word_0/ca
      -- CP-element group 176: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_Update/LOAD_one_475_Merge/$entry
      -- CP-element group 176: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_Update/LOAD_one_475_Merge/$exit
      -- CP-element group 176: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_Update/LOAD_one_475_Merge/merge_req
      -- CP-element group 176: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_one_475_Update/LOAD_one_475_Merge/merge_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(176)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(176)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(176) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_one_475_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_one_475_load_0_ack_1, ack => try1_CP_1680_elements(176)); -- 
    -- CP-element group 177:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	171 
    -- CP-element group 177: successors 
    -- CP-element group 177: marked-successors 
    -- CP-element group 177: 	168 
    -- CP-element group 177: 	171 
    -- CP-element group 177: 	174 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/CONCAT_u1_u32_477_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/CONCAT_u1_u32_477_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/CONCAT_u1_u32_477_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(177)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(177)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(177) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:CONCAT_u1_u32_477_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u1_u32_477_inst_ack_0, ack => try1_CP_1680_elements(177)); -- 
    -- CP-element group 178:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	172 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	183 
    -- CP-element group 178: marked-successors 
    -- CP-element group 178: 	172 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/CONCAT_u1_u32_477_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/CONCAT_u1_u32_477_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/CONCAT_u1_u32_477_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(178)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(178)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(178) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:CONCAT_u1_u32_477_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u1_u32_477_inst_ack_1, ack => try1_CP_1680_elements(178)); -- 
    -- CP-element group 179:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	166 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	181 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	181 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_481_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_481_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_481_Sample/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(179)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(179)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(179) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_NGG_420_delayed_4_0_479_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_2540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(179), ack => W_NGG_420_delayed_4_0_479_inst_req_0); -- 
    try1_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(166) & try1_CP_1680_elements(181);
      gj_try1_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: marked-predecessors 
    -- CP-element group 180: 	182 
    -- CP-element group 180: 	185 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	182 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_481_update_start_
      -- CP-element group 180: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_481_Update/$entry
      -- CP-element group 180: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_481_Update/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(180)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(180)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(180) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_NGG_420_delayed_4_0_479_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_2545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(180), ack => W_NGG_420_delayed_4_0_479_inst_req_1); -- 
    try1_cp_element_group_180: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_180"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(182) & try1_CP_1680_elements(185);
      gj_try1_cp_element_group_180 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 181:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	179 
    -- CP-element group 181: successors 
    -- CP-element group 181: marked-successors 
    -- CP-element group 181: 	164 
    -- CP-element group 181: 	179 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_481_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_481_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_481_Sample/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(181)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(181)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(181) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_NGG_420_delayed_4_0_479_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_NGG_420_delayed_4_0_479_inst_ack_0, ack => try1_CP_1680_elements(181)); -- 
    -- CP-element group 182:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	180 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182: marked-successors 
    -- CP-element group 182: 	180 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_481_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_481_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_481_Update/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(182)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(182)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(182) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_NGG_420_delayed_4_0_479_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_NGG_420_delayed_4_0_479_inst_ack_1, ack => try1_CP_1680_elements(182)); -- 
    -- CP-element group 183:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: 	178 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	185 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u32_u32_485_sample_start_
      -- CP-element group 183: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u32_u32_485_Sample/$entry
      -- CP-element group 183: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u32_u32_485_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(183)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(183)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(183) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u32_u32_485_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(183), ack => ADD_u32_u32_485_inst_req_0); -- 
    try1_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(182) & try1_CP_1680_elements(178) & try1_CP_1680_elements(185);
      gj_try1_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: marked-predecessors 
    -- CP-element group 184: 	186 
    -- CP-element group 184: 	189 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	186 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u32_u32_485_update_start_
      -- CP-element group 184: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u32_u32_485_Update/$entry
      -- CP-element group 184: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u32_u32_485_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(184)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(184)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(184) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u32_u32_485_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(184), ack => ADD_u32_u32_485_inst_req_1); -- 
    try1_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(186) & try1_CP_1680_elements(189);
      gj_try1_cp_element_group_184 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: marked-successors 
    -- CP-element group 185: 	180 
    -- CP-element group 185: 	183 
    -- CP-element group 185: 	172 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u32_u32_485_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u32_u32_485_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u32_u32_485_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(185)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(185)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(185) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u32_u32_485_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_485_inst_ack_0, ack => try1_CP_1680_elements(185)); -- 
    -- CP-element group 186:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186: marked-successors 
    -- CP-element group 186: 	184 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u32_u32_485_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u32_u32_485_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u32_u32_485_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(186)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(186)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(186) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u32_u32_485_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_485_inst_ack_1, ack => try1_CP_1680_elements(186)); -- 
    -- CP-element group 187:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: marked-predecessors 
    -- CP-element group 187: 	189 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	189 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/call_stmt_490_sample_start_
      -- CP-element group 187: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/call_stmt_490_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/call_stmt_490_Sample/crr
      -- 
    -- logger for CP element group try1_CP_1680_elements(187)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(187)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(187) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:call_stmt_490_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_2568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(187), ack => call_stmt_490_call_req_0); -- 
    try1_cp_element_group_187: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_187"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(186) & try1_CP_1680_elements(189);
      gj_try1_cp_element_group_187 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(187), clk => clk, reset => reset); --
    end block;
    -- CP-element group 188:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: marked-predecessors 
    -- CP-element group 188: 	197 
    -- CP-element group 188: 	190 
    -- CP-element group 188: 	193 
    -- CP-element group 188: 	225 
    -- CP-element group 188: 	229 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	190 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/call_stmt_490_update_start_
      -- CP-element group 188: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/call_stmt_490_Update/$entry
      -- CP-element group 188: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/call_stmt_490_Update/ccr
      -- 
    -- logger for CP element group try1_CP_1680_elements(188)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(188)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(188) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:call_stmt_490_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_2573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(188), ack => call_stmt_490_call_req_1); -- 
    try1_cp_element_group_188: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_188"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= try1_CP_1680_elements(197) & try1_CP_1680_elements(190) & try1_CP_1680_elements(193) & try1_CP_1680_elements(225) & try1_CP_1680_elements(229);
      gj_try1_cp_element_group_188 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(188), clk => clk, reset => reset); --
    end block;
    -- CP-element group 189:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	187 
    -- CP-element group 189: successors 
    -- CP-element group 189: marked-successors 
    -- CP-element group 189: 	184 
    -- CP-element group 189: 	187 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/call_stmt_490_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/call_stmt_490_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/call_stmt_490_Sample/cra
      -- 
    -- logger for CP element group try1_CP_1680_elements(189)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(189)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(189) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:call_stmt_490_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_2569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_490_call_ack_0, ack => try1_CP_1680_elements(189)); -- 
    -- CP-element group 190:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	188 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	195 
    -- CP-element group 190: 	191 
    -- CP-element group 190: 	223 
    -- CP-element group 190: 	227 
    -- CP-element group 190: marked-successors 
    -- CP-element group 190: 	188 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/call_stmt_490_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/call_stmt_490_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/call_stmt_490_Update/cca
      -- 
    -- logger for CP element group try1_CP_1680_elements(190)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(190)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(190) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:call_stmt_490_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_2574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_490_call_ack_1, ack => try1_CP_1680_elements(190)); -- 
    -- CP-element group 191:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: marked-predecessors 
    -- CP-element group 191: 	193 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	193 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_493_sample_start_
      -- CP-element group 191: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_493_Sample/$entry
      -- CP-element group 191: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_493_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(191)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(191)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(191) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_493_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(191), ack => slice_493_inst_req_0); -- 
    try1_cp_element_group_191: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_191"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(190) & try1_CP_1680_elements(193);
      gj_try1_cp_element_group_191 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(191), clk => clk, reset => reset); --
    end block;
    -- CP-element group 192:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: marked-predecessors 
    -- CP-element group 192: 	194 
    -- CP-element group 192: 	221 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	194 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_493_update_start_
      -- CP-element group 192: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_493_Update/$entry
      -- CP-element group 192: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_493_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(192)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(192)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(192) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_493_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(192), ack => slice_493_inst_req_1); -- 
    try1_cp_element_group_192: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_192"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(194) & try1_CP_1680_elements(221);
      gj_try1_cp_element_group_192 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(192), clk => clk, reset => reset); --
    end block;
    -- CP-element group 193:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	191 
    -- CP-element group 193: successors 
    -- CP-element group 193: marked-successors 
    -- CP-element group 193: 	188 
    -- CP-element group 193: 	191 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_493_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_493_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_493_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(193)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(193)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(193) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_493_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_493_inst_ack_0, ack => try1_CP_1680_elements(193)); -- 
    -- CP-element group 194:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	192 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	219 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	192 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_493_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_493_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_493_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(194)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(194)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(194) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_493_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_493_inst_ack_1, ack => try1_CP_1680_elements(194)); -- 
    -- CP-element group 195:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	190 
    -- CP-element group 195: marked-predecessors 
    -- CP-element group 195: 	197 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	197 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_497_sample_start_
      -- CP-element group 195: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_497_Sample/$entry
      -- CP-element group 195: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_497_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(195)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(195)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(195) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_497_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(195), ack => slice_497_inst_req_0); -- 
    try1_cp_element_group_195: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_195"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(190) & try1_CP_1680_elements(197);
      gj_try1_cp_element_group_195 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(195), clk => clk, reset => reset); --
    end block;
    -- CP-element group 196:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: marked-predecessors 
    -- CP-element group 196: 	198 
    -- CP-element group 196: 	213 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_497_update_start_
      -- CP-element group 196: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_497_Update/$entry
      -- CP-element group 196: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_497_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(196)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(196)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(196) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_497_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(196), ack => slice_497_inst_req_1); -- 
    try1_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(198) & try1_CP_1680_elements(213);
      gj_try1_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	195 
    -- CP-element group 197: successors 
    -- CP-element group 197: marked-successors 
    -- CP-element group 197: 	195 
    -- CP-element group 197: 	188 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_497_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_497_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_497_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(197)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(197)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(197) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_497_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_497_inst_ack_0, ack => try1_CP_1680_elements(197)); -- 
    -- CP-element group 198:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	211 
    -- CP-element group 198: marked-successors 
    -- CP-element group 198: 	196 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_497_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_497_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_497_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(198)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(198)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(198) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_497_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_497_inst_ack_1, ack => try1_CP_1680_elements(198)); -- 
    -- CP-element group 199:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	204 
    -- CP-element group 199: marked-predecessors 
    -- CP-element group 199: 	205 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	205 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_502_sample_start_
      -- CP-element group 199: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_502_Sample/$entry
      -- CP-element group 199: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_502_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(199)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(199)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(199) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u16_u16_502_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(199), ack => ADD_u16_u16_502_inst_req_0); -- 
    try1_cp_element_group_199: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_199"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(204) & try1_CP_1680_elements(205);
      gj_try1_cp_element_group_199 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(199), clk => clk, reset => reset); --
    end block;
    -- CP-element group 200:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: marked-predecessors 
    -- CP-element group 200: 	217 
    -- CP-element group 200: 	206 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	206 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_502_update_start_
      -- CP-element group 200: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_502_Update/$entry
      -- CP-element group 200: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_502_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(200)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(200)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(200) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u16_u16_502_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(200), ack => ADD_u16_u16_502_inst_req_1); -- 
    try1_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(217) & try1_CP_1680_elements(206);
      gj_try1_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	139 
    -- CP-element group 201: marked-predecessors 
    -- CP-element group 201: 	203 
    -- CP-element group 201: 	277 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	203 
    -- CP-element group 201:  members (5) 
      -- CP-element group 201: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_sample_start_
      -- CP-element group 201: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_Sample/$entry
      -- CP-element group 201: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_Sample/word_access_start/$entry
      -- CP-element group 201: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_Sample/word_access_start/word_0/$entry
      -- CP-element group 201: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(201)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(201)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(201) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_PJ_500_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(201), ack => LOAD_PJ_500_load_0_req_0); -- 
    try1_cp_element_group_201: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_201"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(139) & try1_CP_1680_elements(203) & try1_CP_1680_elements(277);
      gj_try1_cp_element_group_201 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(201), clk => clk, reset => reset); --
    end block;
    -- CP-element group 202:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: marked-predecessors 
    -- CP-element group 202: 	204 
    -- CP-element group 202: 	205 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202:  members (5) 
      -- CP-element group 202: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_update_start_
      -- CP-element group 202: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_Update/$entry
      -- CP-element group 202: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_Update/word_access_complete/$entry
      -- CP-element group 202: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_Update/word_access_complete/word_0/$entry
      -- CP-element group 202: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(202)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(202)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(202) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_PJ_500_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(202), ack => LOAD_PJ_500_load_0_req_1); -- 
    try1_cp_element_group_202: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_202"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(204) & try1_CP_1680_elements(205);
      gj_try1_cp_element_group_202 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(202), clk => clk, reset => reset); --
    end block;
    -- CP-element group 203:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	201 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	283 
    -- CP-element group 203: marked-successors 
    -- CP-element group 203: 	201 
    -- CP-element group 203:  members (5) 
      -- CP-element group 203: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_Sample/word_access_start/$exit
      -- CP-element group 203: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_Sample/word_access_start/word_0/$exit
      -- CP-element group 203: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(203)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(203)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(203) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_PJ_500_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_PJ_500_load_0_ack_0, ack => try1_CP_1680_elements(203)); -- 
    -- CP-element group 204:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	202 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	199 
    -- CP-element group 204: marked-successors 
    -- CP-element group 204: 	202 
    -- CP-element group 204:  members (9) 
      -- CP-element group 204: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_Update/word_access_complete/$exit
      -- CP-element group 204: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_Update/word_access_complete/word_0/$exit
      -- CP-element group 204: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_Update/word_access_complete/word_0/ca
      -- CP-element group 204: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_Update/LOAD_PJ_500_Merge/$entry
      -- CP-element group 204: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_Update/LOAD_PJ_500_Merge/$exit
      -- CP-element group 204: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_Update/LOAD_PJ_500_Merge/merge_req
      -- CP-element group 204: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_Update/LOAD_PJ_500_Merge/merge_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(204)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(204)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(204) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_PJ_500_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_PJ_500_load_0_ack_1, ack => try1_CP_1680_elements(204)); -- 
    -- CP-element group 205:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	199 
    -- CP-element group 205: successors 
    -- CP-element group 205: marked-successors 
    -- CP-element group 205: 	199 
    -- CP-element group 205: 	202 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_502_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_502_Sample/$exit
      -- CP-element group 205: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_502_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(205)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(205)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(205) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u16_u16_502_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_502_inst_ack_0, ack => try1_CP_1680_elements(205)); -- 
    -- CP-element group 206:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	200 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	215 
    -- CP-element group 206: marked-successors 
    -- CP-element group 206: 	200 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_502_update_completed_
      -- CP-element group 206: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_502_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_502_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(206)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(206)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(206) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u16_u16_502_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_502_inst_ack_1, ack => try1_CP_1680_elements(206)); -- 
    -- CP-element group 207:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	139 
    -- CP-element group 207: marked-predecessors 
    -- CP-element group 207: 	277 
    -- CP-element group 207: 	209 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	209 
    -- CP-element group 207:  members (5) 
      -- CP-element group 207: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_Sample/word_access_start/$entry
      -- CP-element group 207: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_Sample/word_access_start/word_0/$entry
      -- CP-element group 207: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(207)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(207)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(207) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_PJ_505_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(207), ack => LOAD_PJ_505_load_0_req_0); -- 
    try1_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(139) & try1_CP_1680_elements(277) & try1_CP_1680_elements(209);
      gj_try1_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: marked-predecessors 
    -- CP-element group 208: 	213 
    -- CP-element group 208: 	210 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (5) 
      -- CP-element group 208: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_update_start_
      -- CP-element group 208: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_Update/word_access_complete/$entry
      -- CP-element group 208: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_Update/word_access_complete/word_0/$entry
      -- CP-element group 208: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(208)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(208)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(208) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_PJ_505_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(208), ack => LOAD_PJ_505_load_0_req_1); -- 
    try1_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(213) & try1_CP_1680_elements(210);
      gj_try1_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	207 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	284 
    -- CP-element group 209: marked-successors 
    -- CP-element group 209: 	207 
    -- CP-element group 209:  members (5) 
      -- CP-element group 209: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_sample_completed_
      -- CP-element group 209: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_Sample/$exit
      -- CP-element group 209: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_Sample/word_access_start/$exit
      -- CP-element group 209: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_Sample/word_access_start/word_0/$exit
      -- CP-element group 209: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(209)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(209)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(209) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_PJ_505_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_PJ_505_load_0_ack_0, ack => try1_CP_1680_elements(209)); -- 
    -- CP-element group 210:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210: marked-successors 
    -- CP-element group 210: 	208 
    -- CP-element group 210:  members (35) 
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_update_completed_
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_Update/$exit
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_Update/word_access_complete/$exit
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_Update/word_access_complete/word_0/$exit
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_Update/word_access_complete/word_0/ca
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_Update/LOAD_PJ_505_Merge/$entry
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_Update/LOAD_PJ_505_Merge/$exit
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_Update/LOAD_PJ_505_Merge/merge_req
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_Update/LOAD_PJ_505_Merge/merge_ack
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_word_address_calculated
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_root_address_calculated
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_offset_calculated
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_index_resized_0
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_index_scaled_0
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_index_computed_0
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_index_resize_0/$entry
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_index_resize_0/$exit
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_index_resize_0/index_resize_req
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_index_resize_0/index_resize_ack
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_index_scale_0/$entry
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_index_scale_0/$exit
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_index_scale_0/scale_rename_req
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_index_scale_0/scale_rename_ack
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_final_index_sum_regn/$entry
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_final_index_sum_regn/$exit
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_final_index_sum_regn/req
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_final_index_sum_regn/ack
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_base_plus_offset/$entry
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_base_plus_offset/$exit
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_base_plus_offset/sum_rename_req
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_base_plus_offset/sum_rename_ack
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_word_addrgen/$entry
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_word_addrgen/$exit
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_word_addrgen/root_register_req
      -- CP-element group 210: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(210)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(210)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(210) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_PJ_505_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_PJ_505_load_0_ack_1, ack => try1_CP_1680_elements(210)); -- 
    -- CP-element group 211:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	198 
    -- CP-element group 211: 	210 
    -- CP-element group 211: marked-predecessors 
    -- CP-element group 211: 	261 
    -- CP-element group 211: 	213 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (9) 
      -- CP-element group 211: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_sample_start_
      -- CP-element group 211: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_Sample/$entry
      -- CP-element group 211: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_Sample/array_obj_ref_508_Split/$entry
      -- CP-element group 211: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_Sample/array_obj_ref_508_Split/$exit
      -- CP-element group 211: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_Sample/array_obj_ref_508_Split/split_req
      -- CP-element group 211: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_Sample/array_obj_ref_508_Split/split_ack
      -- CP-element group 211: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_Sample/word_access_start/$entry
      -- CP-element group 211: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_Sample/word_access_start/word_0/$entry
      -- CP-element group 211: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(211)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(211)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(211) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_508_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(211), ack => array_obj_ref_508_store_0_req_0); -- 
    try1_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= try1_CP_1680_elements(198) & try1_CP_1680_elements(210) & try1_CP_1680_elements(261) & try1_CP_1680_elements(213);
      gj_try1_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: marked-predecessors 
    -- CP-element group 212: 	214 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	214 
    -- CP-element group 212:  members (5) 
      -- CP-element group 212: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_update_start_
      -- CP-element group 212: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_Update/$entry
      -- CP-element group 212: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_Update/word_access_complete/$entry
      -- CP-element group 212: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_Update/word_access_complete/word_0/$entry
      -- CP-element group 212: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(212)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(212)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(212) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_508_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(212), ack => array_obj_ref_508_store_0_req_1); -- 
    try1_cp_element_group_212: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_212"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(214);
      gj_try1_cp_element_group_212 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(212), clk => clk, reset => reset); --
    end block;
    -- CP-element group 213:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	280 
    -- CP-element group 213: marked-successors 
    -- CP-element group 213: 	196 
    -- CP-element group 213: 	208 
    -- CP-element group 213: 	211 
    -- CP-element group 213:  members (5) 
      -- CP-element group 213: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_Sample/word_access_start/$exit
      -- CP-element group 213: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_Sample/word_access_start/word_0/$exit
      -- CP-element group 213: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(213)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(213)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(213) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_508_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_508_store_0_ack_0, ack => try1_CP_1680_elements(213)); -- 
    -- CP-element group 214:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	212 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	288 
    -- CP-element group 214: marked-successors 
    -- CP-element group 214: 	212 
    -- CP-element group 214:  members (5) 
      -- CP-element group 214: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_Update/word_access_complete/$exit
      -- CP-element group 214: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_Update/word_access_complete/word_0/$exit
      -- CP-element group 214: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(214)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(214)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(214) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_508_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_508_store_0_ack_1, ack => try1_CP_1680_elements(214)); -- 
    -- CP-element group 215:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	206 
    -- CP-element group 215: marked-predecessors 
    -- CP-element group 215: 	217 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	217 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_513_sample_start_
      -- CP-element group 215: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_513_Sample/$entry
      -- CP-element group 215: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_513_Sample/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(215)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(215)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(215) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_PPJ_444_delayed_6_0_511_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_2752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(215), ack => W_PPJ_444_delayed_6_0_511_inst_req_0); -- 
    try1_cp_element_group_215: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_215"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(206) & try1_CP_1680_elements(217);
      gj_try1_cp_element_group_215 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(215), clk => clk, reset => reset); --
    end block;
    -- CP-element group 216:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: marked-predecessors 
    -- CP-element group 216: 	218 
    -- CP-element group 216: 	221 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	218 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_513_update_start_
      -- CP-element group 216: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_513_Update/$entry
      -- CP-element group 216: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_513_Update/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(216)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(216)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(216) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_PPJ_444_delayed_6_0_511_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_2757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(216), ack => W_PPJ_444_delayed_6_0_511_inst_req_1); -- 
    try1_cp_element_group_216: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_216"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(218) & try1_CP_1680_elements(221);
      gj_try1_cp_element_group_216 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(216), clk => clk, reset => reset); --
    end block;
    -- CP-element group 217:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	215 
    -- CP-element group 217: successors 
    -- CP-element group 217: marked-successors 
    -- CP-element group 217: 	200 
    -- CP-element group 217: 	215 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_513_sample_completed_
      -- CP-element group 217: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_513_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_513_Sample/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(217)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(217)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(217) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_PPJ_444_delayed_6_0_511_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_PPJ_444_delayed_6_0_511_inst_ack_0, ack => try1_CP_1680_elements(217)); -- 
    -- CP-element group 218:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	216 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218: marked-successors 
    -- CP-element group 218: 	216 
    -- CP-element group 218:  members (29) 
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_513_update_completed_
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_513_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_513_Update/ack
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_word_address_calculated
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_root_address_calculated
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_offset_calculated
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_index_resized_0
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_index_scaled_0
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_index_computed_0
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_index_resize_0/$entry
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_index_resize_0/$exit
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_index_resize_0/index_resize_req
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_index_resize_0/index_resize_ack
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_index_scale_0/$entry
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_index_scale_0/$exit
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_index_scale_0/scale_rename_req
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_index_scale_0/scale_rename_ack
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_final_index_sum_regn/$entry
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_final_index_sum_regn/$exit
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_final_index_sum_regn/req
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_final_index_sum_regn/ack
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_base_plus_offset/$entry
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_base_plus_offset/$exit
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_base_plus_offset/sum_rename_req
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_base_plus_offset/sum_rename_ack
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_word_addrgen/$entry
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_word_addrgen/$exit
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_word_addrgen/root_register_req
      -- CP-element group 218: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(218)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(218)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(218) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_PPJ_444_delayed_6_0_511_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_PPJ_444_delayed_6_0_511_inst_ack_1, ack => try1_CP_1680_elements(218)); -- 
    -- CP-element group 219:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	194 
    -- CP-element group 219: 	218 
    -- CP-element group 219: 	280 
    -- CP-element group 219: marked-predecessors 
    -- CP-element group 219: 	221 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (9) 
      -- CP-element group 219: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_sample_start_
      -- CP-element group 219: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_Sample/$entry
      -- CP-element group 219: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_Sample/array_obj_ref_515_Split/$entry
      -- CP-element group 219: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_Sample/array_obj_ref_515_Split/$exit
      -- CP-element group 219: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_Sample/array_obj_ref_515_Split/split_req
      -- CP-element group 219: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_Sample/array_obj_ref_515_Split/split_ack
      -- CP-element group 219: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_Sample/word_access_start/$entry
      -- CP-element group 219: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_Sample/word_access_start/word_0/$entry
      -- CP-element group 219: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(219)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(219)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(219) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_515_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(219), ack => array_obj_ref_515_store_0_req_0); -- 
    try1_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= try1_CP_1680_elements(194) & try1_CP_1680_elements(218) & try1_CP_1680_elements(280) & try1_CP_1680_elements(221);
      gj_try1_cp_element_group_219 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: marked-predecessors 
    -- CP-element group 220: 	222 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	222 
    -- CP-element group 220:  members (5) 
      -- CP-element group 220: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_update_start_
      -- CP-element group 220: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_Update/$entry
      -- CP-element group 220: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_Update/word_access_complete/$entry
      -- CP-element group 220: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_Update/word_access_complete/word_0/$entry
      -- CP-element group 220: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(220)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(220)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(220) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_515_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(220), ack => array_obj_ref_515_store_0_req_1); -- 
    try1_cp_element_group_220: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_220"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(222);
      gj_try1_cp_element_group_220 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(220), clk => clk, reset => reset); --
    end block;
    -- CP-element group 221:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	281 
    -- CP-element group 221: marked-successors 
    -- CP-element group 221: 	192 
    -- CP-element group 221: 	216 
    -- CP-element group 221: 	219 
    -- CP-element group 221:  members (5) 
      -- CP-element group 221: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_sample_completed_
      -- CP-element group 221: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_Sample/$exit
      -- CP-element group 221: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_Sample/word_access_start/$exit
      -- CP-element group 221: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_Sample/word_access_start/word_0/$exit
      -- CP-element group 221: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(221)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(221)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(221) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_515_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_515_store_0_ack_0, ack => try1_CP_1680_elements(221)); -- 
    -- CP-element group 222:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	220 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	288 
    -- CP-element group 222: marked-successors 
    -- CP-element group 222: 	220 
    -- CP-element group 222:  members (5) 
      -- CP-element group 222: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_update_completed_
      -- CP-element group 222: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_Update/word_access_complete/$exit
      -- CP-element group 222: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_Update/word_access_complete/word_0/$exit
      -- CP-element group 222: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(222)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(222)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(222) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_515_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_515_store_0_ack_1, ack => try1_CP_1680_elements(222)); -- 
    -- CP-element group 223:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	190 
    -- CP-element group 223: marked-predecessors 
    -- CP-element group 223: 	225 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	225 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_520_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_520_Sample/$entry
      -- CP-element group 223: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_520_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(223)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(223)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(223) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_520_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(223), ack => slice_520_inst_req_0); -- 
    try1_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(190) & try1_CP_1680_elements(225);
      gj_try1_cp_element_group_223 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: marked-predecessors 
    -- CP-element group 224: 	261 
    -- CP-element group 224: 	226 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	226 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_520_update_start_
      -- CP-element group 224: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_520_Update/$entry
      -- CP-element group 224: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_520_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(224)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(224)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(224) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_520_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(224), ack => slice_520_inst_req_1); -- 
    try1_cp_element_group_224: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_224"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(261) & try1_CP_1680_elements(226);
      gj_try1_cp_element_group_224 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(224), clk => clk, reset => reset); --
    end block;
    -- CP-element group 225:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	223 
    -- CP-element group 225: successors 
    -- CP-element group 225: marked-successors 
    -- CP-element group 225: 	188 
    -- CP-element group 225: 	223 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_520_sample_completed_
      -- CP-element group 225: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_520_Sample/$exit
      -- CP-element group 225: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_520_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(225)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(225)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(225) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_520_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_520_inst_ack_0, ack => try1_CP_1680_elements(225)); -- 
    -- CP-element group 226:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	224 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	259 
    -- CP-element group 226: marked-successors 
    -- CP-element group 226: 	224 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_520_update_completed_
      -- CP-element group 226: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_520_Update/$exit
      -- CP-element group 226: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_520_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(226)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(226)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(226) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_520_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_520_inst_ack_1, ack => try1_CP_1680_elements(226)); -- 
    -- CP-element group 227:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	190 
    -- CP-element group 227: marked-predecessors 
    -- CP-element group 227: 	229 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	229 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_524_sample_start_
      -- CP-element group 227: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_524_Sample/$entry
      -- CP-element group 227: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_524_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(227)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(227)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(227) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_524_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(227), ack => slice_524_inst_req_0); -- 
    try1_cp_element_group_227: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_227"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(190) & try1_CP_1680_elements(229);
      gj_try1_cp_element_group_227 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(227), clk => clk, reset => reset); --
    end block;
    -- CP-element group 228:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: marked-predecessors 
    -- CP-element group 228: 	253 
    -- CP-element group 228: 	230 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_524_update_start_
      -- CP-element group 228: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_524_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_524_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(228)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(228)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(228) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_524_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(228), ack => slice_524_inst_req_1); -- 
    try1_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(253) & try1_CP_1680_elements(230);
      gj_try1_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	227 
    -- CP-element group 229: successors 
    -- CP-element group 229: marked-successors 
    -- CP-element group 229: 	188 
    -- CP-element group 229: 	227 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_524_sample_completed_
      -- CP-element group 229: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_524_Sample/$exit
      -- CP-element group 229: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_524_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(229)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(229)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(229) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_524_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_524_inst_ack_0, ack => try1_CP_1680_elements(229)); -- 
    -- CP-element group 230:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	251 
    -- CP-element group 230: marked-successors 
    -- CP-element group 230: 	228 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_524_update_completed_
      -- CP-element group 230: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_524_Update/$exit
      -- CP-element group 230: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/slice_524_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(230)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(230)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(230) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_524_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_524_inst_ack_1, ack => try1_CP_1680_elements(230)); -- 
    -- CP-element group 231:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	236 
    -- CP-element group 231: marked-predecessors 
    -- CP-element group 231: 	237 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	237 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_529_sample_start_
      -- CP-element group 231: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_529_Sample/$entry
      -- CP-element group 231: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_529_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(231)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(231)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(231) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u16_u16_529_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(231), ack => ADD_u16_u16_529_inst_req_0); -- 
    try1_cp_element_group_231: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_231"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(236) & try1_CP_1680_elements(237);
      gj_try1_cp_element_group_231 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(231), clk => clk, reset => reset); --
    end block;
    -- CP-element group 232:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: marked-predecessors 
    -- CP-element group 232: 	238 
    -- CP-element group 232: 	249 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	238 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_529_update_start_
      -- CP-element group 232: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_529_Update/$entry
      -- CP-element group 232: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_529_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(232)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(232)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(232) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u16_u16_529_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(232), ack => ADD_u16_u16_529_inst_req_1); -- 
    try1_cp_element_group_232: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_232"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(238) & try1_CP_1680_elements(249);
      gj_try1_cp_element_group_232 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(232), clk => clk, reset => reset); --
    end block;
    -- CP-element group 233:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	139 
    -- CP-element group 233: marked-predecessors 
    -- CP-element group 233: 	277 
    -- CP-element group 233: 	235 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	235 
    -- CP-element group 233:  members (5) 
      -- CP-element group 233: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_sample_start_
      -- CP-element group 233: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_Sample/$entry
      -- CP-element group 233: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_Sample/word_access_start/$entry
      -- CP-element group 233: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_Sample/word_access_start/word_0/$entry
      -- CP-element group 233: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(233)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(233)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(233) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_PJ_527_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(233), ack => LOAD_PJ_527_load_0_req_0); -- 
    try1_cp_element_group_233: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_233"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(139) & try1_CP_1680_elements(277) & try1_CP_1680_elements(235);
      gj_try1_cp_element_group_233 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(233), clk => clk, reset => reset); --
    end block;
    -- CP-element group 234:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: marked-predecessors 
    -- CP-element group 234: 	236 
    -- CP-element group 234: 	237 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (5) 
      -- CP-element group 234: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_update_start_
      -- CP-element group 234: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_Update/word_access_complete/$entry
      -- CP-element group 234: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_Update/word_access_complete/word_0/$entry
      -- CP-element group 234: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(234)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(234)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(234) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_PJ_527_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(234), ack => LOAD_PJ_527_load_0_req_1); -- 
    try1_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(236) & try1_CP_1680_elements(237);
      gj_try1_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	233 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	285 
    -- CP-element group 235: marked-successors 
    -- CP-element group 235: 	233 
    -- CP-element group 235:  members (5) 
      -- CP-element group 235: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_Sample/word_access_start/$exit
      -- CP-element group 235: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_Sample/word_access_start/word_0/$exit
      -- CP-element group 235: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(235)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(235)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(235) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_PJ_527_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_PJ_527_load_0_ack_0, ack => try1_CP_1680_elements(235)); -- 
    -- CP-element group 236:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	231 
    -- CP-element group 236: marked-successors 
    -- CP-element group 236: 	234 
    -- CP-element group 236:  members (9) 
      -- CP-element group 236: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_Update/word_access_complete/$exit
      -- CP-element group 236: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_Update/word_access_complete/word_0/$exit
      -- CP-element group 236: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_Update/word_access_complete/word_0/ca
      -- CP-element group 236: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_Update/LOAD_PJ_527_Merge/$entry
      -- CP-element group 236: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_Update/LOAD_PJ_527_Merge/$exit
      -- CP-element group 236: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_Update/LOAD_PJ_527_Merge/merge_req
      -- CP-element group 236: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_Update/LOAD_PJ_527_Merge/merge_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(236)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(236)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(236) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_PJ_527_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_PJ_527_load_0_ack_1, ack => try1_CP_1680_elements(236)); -- 
    -- CP-element group 237:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	231 
    -- CP-element group 237: successors 
    -- CP-element group 237: marked-successors 
    -- CP-element group 237: 	231 
    -- CP-element group 237: 	234 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_529_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_529_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_529_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(237)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(237)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(237) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u16_u16_529_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_529_inst_ack_0, ack => try1_CP_1680_elements(237)); -- 
    -- CP-element group 238:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	232 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	247 
    -- CP-element group 238: marked-successors 
    -- CP-element group 238: 	232 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_529_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_529_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_529_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(238)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(238)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(238) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u16_u16_529_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_529_inst_ack_1, ack => try1_CP_1680_elements(238)); -- 
    -- CP-element group 239:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	244 
    -- CP-element group 239: marked-predecessors 
    -- CP-element group 239: 	245 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	245 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_534_sample_start_
      -- CP-element group 239: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_534_Sample/$entry
      -- CP-element group 239: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_534_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(239)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(239)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(239) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u16_u16_534_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(239), ack => ADD_u16_u16_534_inst_req_0); -- 
    try1_cp_element_group_239: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_239"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(244) & try1_CP_1680_elements(245);
      gj_try1_cp_element_group_239 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(239), clk => clk, reset => reset); --
    end block;
    -- CP-element group 240:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: marked-predecessors 
    -- CP-element group 240: 	257 
    -- CP-element group 240: 	246 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	246 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_534_update_start_
      -- CP-element group 240: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_534_Update/$entry
      -- CP-element group 240: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_534_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(240)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(240)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(240) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u16_u16_534_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(240), ack => ADD_u16_u16_534_inst_req_1); -- 
    try1_cp_element_group_240: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_240"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(257) & try1_CP_1680_elements(246);
      gj_try1_cp_element_group_240 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(240), clk => clk, reset => reset); --
    end block;
    -- CP-element group 241:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	139 
    -- CP-element group 241: marked-predecessors 
    -- CP-element group 241: 	277 
    -- CP-element group 241: 	243 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	243 
    -- CP-element group 241:  members (5) 
      -- CP-element group 241: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_sample_start_
      -- CP-element group 241: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_Sample/$entry
      -- CP-element group 241: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_Sample/word_access_start/$entry
      -- CP-element group 241: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_Sample/word_access_start/word_0/$entry
      -- CP-element group 241: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(241)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(241)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(241) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_PJ_532_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(241), ack => LOAD_PJ_532_load_0_req_0); -- 
    try1_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(139) & try1_CP_1680_elements(277) & try1_CP_1680_elements(243);
      gj_try1_cp_element_group_241 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: marked-predecessors 
    -- CP-element group 242: 	244 
    -- CP-element group 242: 	245 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (5) 
      -- CP-element group 242: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_update_start_
      -- CP-element group 242: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_Update/$entry
      -- CP-element group 242: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_Update/word_access_complete/$entry
      -- CP-element group 242: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_Update/word_access_complete/word_0/$entry
      -- CP-element group 242: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(242)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(242)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(242) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_PJ_532_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(242), ack => LOAD_PJ_532_load_0_req_1); -- 
    try1_cp_element_group_242: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_242"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(244) & try1_CP_1680_elements(245);
      gj_try1_cp_element_group_242 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(242), clk => clk, reset => reset); --
    end block;
    -- CP-element group 243:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	241 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	286 
    -- CP-element group 243: marked-successors 
    -- CP-element group 243: 	241 
    -- CP-element group 243:  members (5) 
      -- CP-element group 243: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_Sample/word_access_start/$exit
      -- CP-element group 243: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_Sample/word_access_start/word_0/$exit
      -- CP-element group 243: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(243)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(243)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(243) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_PJ_532_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_PJ_532_load_0_ack_0, ack => try1_CP_1680_elements(243)); -- 
    -- CP-element group 244:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	239 
    -- CP-element group 244: marked-successors 
    -- CP-element group 244: 	242 
    -- CP-element group 244:  members (9) 
      -- CP-element group 244: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_Update/word_access_complete/$exit
      -- CP-element group 244: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_Update/word_access_complete/word_0/$exit
      -- CP-element group 244: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_Update/word_access_complete/word_0/ca
      -- CP-element group 244: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_Update/LOAD_PJ_532_Merge/$entry
      -- CP-element group 244: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_Update/LOAD_PJ_532_Merge/$exit
      -- CP-element group 244: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_Update/LOAD_PJ_532_Merge/merge_req
      -- CP-element group 244: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_Update/LOAD_PJ_532_Merge/merge_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(244)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(244)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(244) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_PJ_532_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_PJ_532_load_0_ack_1, ack => try1_CP_1680_elements(244)); -- 
    -- CP-element group 245:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	239 
    -- CP-element group 245: successors 
    -- CP-element group 245: marked-successors 
    -- CP-element group 245: 	239 
    -- CP-element group 245: 	242 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_534_sample_completed_
      -- CP-element group 245: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_534_Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_534_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(245)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(245)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(245) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u16_u16_534_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_534_inst_ack_0, ack => try1_CP_1680_elements(245)); -- 
    -- CP-element group 246:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	240 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	255 
    -- CP-element group 246: marked-successors 
    -- CP-element group 246: 	240 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_534_update_completed_
      -- CP-element group 246: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_534_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_534_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(246)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(246)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(246) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u16_u16_534_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_534_inst_ack_1, ack => try1_CP_1680_elements(246)); -- 
    -- CP-element group 247:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	238 
    -- CP-element group 247: marked-predecessors 
    -- CP-element group 247: 	249 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	249 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_538_sample_start_
      -- CP-element group 247: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_538_Sample/$entry
      -- CP-element group 247: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_538_Sample/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(247)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(247)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(247) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_PPPJ_466_delayed_6_0_536_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_2950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(247), ack => W_PPPJ_466_delayed_6_0_536_inst_req_0); -- 
    try1_cp_element_group_247: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_247"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(238) & try1_CP_1680_elements(249);
      gj_try1_cp_element_group_247 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(247), clk => clk, reset => reset); --
    end block;
    -- CP-element group 248:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: marked-predecessors 
    -- CP-element group 248: 	253 
    -- CP-element group 248: 	250 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	250 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_538_update_start_
      -- CP-element group 248: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_538_Update/$entry
      -- CP-element group 248: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_538_Update/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(248)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(248)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(248) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_PPPJ_466_delayed_6_0_536_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_2955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(248), ack => W_PPPJ_466_delayed_6_0_536_inst_req_1); -- 
    try1_cp_element_group_248: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_248"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(253) & try1_CP_1680_elements(250);
      gj_try1_cp_element_group_248 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(248), clk => clk, reset => reset); --
    end block;
    -- CP-element group 249:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	247 
    -- CP-element group 249: successors 
    -- CP-element group 249: marked-successors 
    -- CP-element group 249: 	232 
    -- CP-element group 249: 	247 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_538_sample_completed_
      -- CP-element group 249: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_538_Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_538_Sample/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(249)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(249)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(249) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_PPPJ_466_delayed_6_0_536_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_PPPJ_466_delayed_6_0_536_inst_ack_0, ack => try1_CP_1680_elements(249)); -- 
    -- CP-element group 250:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	248 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250: marked-successors 
    -- CP-element group 250: 	248 
    -- CP-element group 250:  members (29) 
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_538_update_completed_
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_538_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_538_Update/ack
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_word_address_calculated
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_root_address_calculated
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_offset_calculated
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_index_resized_0
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_index_scaled_0
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_index_computed_0
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_index_resize_0/$entry
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_index_resize_0/$exit
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_index_resize_0/index_resize_req
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_index_resize_0/index_resize_ack
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_index_scale_0/$entry
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_index_scale_0/$exit
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_index_scale_0/scale_rename_req
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_index_scale_0/scale_rename_ack
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_final_index_sum_regn/$entry
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_final_index_sum_regn/$exit
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_final_index_sum_regn/req
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_final_index_sum_regn/ack
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_base_plus_offset/$entry
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_base_plus_offset/$exit
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_base_plus_offset/sum_rename_req
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_base_plus_offset/sum_rename_ack
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_word_addrgen/$entry
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_word_addrgen/$exit
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_word_addrgen/root_register_req
      -- CP-element group 250: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(250)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(250)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(250) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_PPPJ_466_delayed_6_0_536_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_PPPJ_466_delayed_6_0_536_inst_ack_1, ack => try1_CP_1680_elements(250)); -- 
    -- CP-element group 251:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	281 
    -- CP-element group 251: 	230 
    -- CP-element group 251: 	250 
    -- CP-element group 251: marked-predecessors 
    -- CP-element group 251: 	253 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	253 
    -- CP-element group 251:  members (9) 
      -- CP-element group 251: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_sample_start_
      -- CP-element group 251: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_Sample/$entry
      -- CP-element group 251: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_Sample/array_obj_ref_540_Split/$entry
      -- CP-element group 251: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_Sample/array_obj_ref_540_Split/$exit
      -- CP-element group 251: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_Sample/array_obj_ref_540_Split/split_req
      -- CP-element group 251: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_Sample/array_obj_ref_540_Split/split_ack
      -- CP-element group 251: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_Sample/word_access_start/$entry
      -- CP-element group 251: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_Sample/word_access_start/word_0/$entry
      -- CP-element group 251: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(251)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(251)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(251) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_540_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(251), ack => array_obj_ref_540_store_0_req_0); -- 
    try1_cp_element_group_251: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_251"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= try1_CP_1680_elements(281) & try1_CP_1680_elements(230) & try1_CP_1680_elements(250) & try1_CP_1680_elements(253);
      gj_try1_cp_element_group_251 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(251), clk => clk, reset => reset); --
    end block;
    -- CP-element group 252:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: marked-predecessors 
    -- CP-element group 252: 	254 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	254 
    -- CP-element group 252:  members (5) 
      -- CP-element group 252: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_update_start_
      -- CP-element group 252: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_Update/$entry
      -- CP-element group 252: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_Update/word_access_complete/$entry
      -- CP-element group 252: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_Update/word_access_complete/word_0/$entry
      -- CP-element group 252: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(252)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(252)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(252) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_540_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(252), ack => array_obj_ref_540_store_0_req_1); -- 
    try1_cp_element_group_252: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_252"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(254);
      gj_try1_cp_element_group_252 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(252), clk => clk, reset => reset); --
    end block;
    -- CP-element group 253:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	251 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	282 
    -- CP-element group 253: marked-successors 
    -- CP-element group 253: 	228 
    -- CP-element group 253: 	248 
    -- CP-element group 253: 	251 
    -- CP-element group 253:  members (5) 
      -- CP-element group 253: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_sample_completed_
      -- CP-element group 253: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_Sample/word_access_start/$exit
      -- CP-element group 253: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_Sample/word_access_start/word_0/$exit
      -- CP-element group 253: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(253)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(253)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(253) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_540_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_540_store_0_ack_0, ack => try1_CP_1680_elements(253)); -- 
    -- CP-element group 254:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	252 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	288 
    -- CP-element group 254: marked-successors 
    -- CP-element group 254: 	252 
    -- CP-element group 254:  members (5) 
      -- CP-element group 254: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_update_completed_
      -- CP-element group 254: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_Update/word_access_complete/$exit
      -- CP-element group 254: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_Update/word_access_complete/word_0/$exit
      -- CP-element group 254: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(254)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(254)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(254) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_540_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_540_store_0_ack_1, ack => try1_CP_1680_elements(254)); -- 
    -- CP-element group 255:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	246 
    -- CP-element group 255: marked-predecessors 
    -- CP-element group 255: 	257 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	257 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_545_sample_start_
      -- CP-element group 255: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_545_Sample/$entry
      -- CP-element group 255: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_545_Sample/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(255)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(255)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(255) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_PPPPJ_470_delayed_6_0_543_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(255), ack => W_PPPPJ_470_delayed_6_0_543_inst_req_0); -- 
    try1_cp_element_group_255: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_255"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(246) & try1_CP_1680_elements(257);
      gj_try1_cp_element_group_255 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(255), clk => clk, reset => reset); --
    end block;
    -- CP-element group 256:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: marked-predecessors 
    -- CP-element group 256: 	258 
    -- CP-element group 256: 	261 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	258 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_545_update_start_
      -- CP-element group 256: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_545_Update/$entry
      -- CP-element group 256: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_545_Update/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(256)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(256)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(256) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_PPPPJ_470_delayed_6_0_543_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(256), ack => W_PPPPJ_470_delayed_6_0_543_inst_req_1); -- 
    try1_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(258) & try1_CP_1680_elements(261);
      gj_try1_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	255 
    -- CP-element group 257: successors 
    -- CP-element group 257: marked-successors 
    -- CP-element group 257: 	255 
    -- CP-element group 257: 	240 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_545_sample_completed_
      -- CP-element group 257: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_545_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_545_Sample/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(257)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(257)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(257) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_PPPPJ_470_delayed_6_0_543_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_PPPPJ_470_delayed_6_0_543_inst_ack_0, ack => try1_CP_1680_elements(257)); -- 
    -- CP-element group 258:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	256 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258: marked-successors 
    -- CP-element group 258: 	256 
    -- CP-element group 258:  members (29) 
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_545_update_completed_
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_545_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/assign_stmt_545_Update/ack
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_word_address_calculated
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_root_address_calculated
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_offset_calculated
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_index_resized_0
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_index_scaled_0
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_index_computed_0
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_index_resize_0/$entry
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_index_resize_0/$exit
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_index_resize_0/index_resize_req
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_index_resize_0/index_resize_ack
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_index_scale_0/$entry
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_index_scale_0/$exit
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_index_scale_0/scale_rename_req
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_index_scale_0/scale_rename_ack
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_final_index_sum_regn/$entry
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_final_index_sum_regn/$exit
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_final_index_sum_regn/req
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_final_index_sum_regn/ack
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_base_plus_offset/$entry
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_base_plus_offset/$exit
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_base_plus_offset/sum_rename_req
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_base_plus_offset/sum_rename_ack
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_word_addrgen/$entry
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_word_addrgen/$exit
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_word_addrgen/root_register_req
      -- CP-element group 258: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(258)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(258)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(258) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_PPPPJ_470_delayed_6_0_543_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_PPPPJ_470_delayed_6_0_543_inst_ack_1, ack => try1_CP_1680_elements(258)); -- 
    -- CP-element group 259:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: 	282 
    -- CP-element group 259: 	226 
    -- CP-element group 259: marked-predecessors 
    -- CP-element group 259: 	261 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	261 
    -- CP-element group 259:  members (9) 
      -- CP-element group 259: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_sample_start_
      -- CP-element group 259: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_Sample/$entry
      -- CP-element group 259: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_Sample/array_obj_ref_547_Split/$entry
      -- CP-element group 259: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_Sample/array_obj_ref_547_Split/$exit
      -- CP-element group 259: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_Sample/array_obj_ref_547_Split/split_req
      -- CP-element group 259: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_Sample/array_obj_ref_547_Split/split_ack
      -- CP-element group 259: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_Sample/word_access_start/$entry
      -- CP-element group 259: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_Sample/word_access_start/word_0/$entry
      -- CP-element group 259: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(259)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(259)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(259) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_547_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(259), ack => array_obj_ref_547_store_0_req_0); -- 
    try1_cp_element_group_259: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_259"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= try1_CP_1680_elements(258) & try1_CP_1680_elements(282) & try1_CP_1680_elements(226) & try1_CP_1680_elements(261);
      gj_try1_cp_element_group_259 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(259), clk => clk, reset => reset); --
    end block;
    -- CP-element group 260:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: marked-predecessors 
    -- CP-element group 260: 	262 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	262 
    -- CP-element group 260:  members (5) 
      -- CP-element group 260: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_update_start_
      -- CP-element group 260: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_Update/$entry
      -- CP-element group 260: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_Update/word_access_complete/$entry
      -- CP-element group 260: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_Update/word_access_complete/word_0/$entry
      -- CP-element group 260: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(260)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(260)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(260) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_547_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(260), ack => array_obj_ref_547_store_0_req_1); -- 
    try1_cp_element_group_260: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_260"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(262);
      gj_try1_cp_element_group_260 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(260), clk => clk, reset => reset); --
    end block;
    -- CP-element group 261:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	259 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	288 
    -- CP-element group 261: marked-successors 
    -- CP-element group 261: 	256 
    -- CP-element group 261: 	259 
    -- CP-element group 261: 	211 
    -- CP-element group 261: 	224 
    -- CP-element group 261:  members (6) 
      -- CP-element group 261: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_sample_completed_
      -- CP-element group 261: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_Sample/word_access_start/$exit
      -- CP-element group 261: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_Sample/word_access_start/word_0/$exit
      -- CP-element group 261: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_Sample/word_access_start/word_0/ra
      -- CP-element group 261: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ring_reenable_memory_space_3
      -- 
    -- logger for CP element group try1_CP_1680_elements(261)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(261)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(261) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_547_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_547_store_0_ack_0, ack => try1_CP_1680_elements(261)); -- 
    -- CP-element group 262:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	260 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	288 
    -- CP-element group 262: marked-successors 
    -- CP-element group 262: 	260 
    -- CP-element group 262:  members (5) 
      -- CP-element group 262: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_update_completed_
      -- CP-element group 262: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_Update/word_access_complete/$exit
      -- CP-element group 262: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_Update/word_access_complete/word_0/$exit
      -- CP-element group 262: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_547_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(262)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(262)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(262) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_547_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_547_store_0_ack_1, ack => try1_CP_1680_elements(262)); -- 
    -- CP-element group 263:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	145 
    -- CP-element group 263: marked-predecessors 
    -- CP-element group 263: 	265 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	265 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u12_u12_553_Sample/$entry
      -- CP-element group 263: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u12_u12_553_Sample/rr
      -- CP-element group 263: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u12_u12_553_sample_start_
      -- 
    -- logger for CP element group try1_CP_1680_elements(263)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(263)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(263) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_553_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(263), ack => ADD_u12_u12_553_inst_req_0); -- 
    try1_cp_element_group_263: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_263"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(145) & try1_CP_1680_elements(265);
      gj_try1_cp_element_group_263 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(263), clk => clk, reset => reset); --
    end block;
    -- CP-element group 264:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	144 
    -- CP-element group 264: marked-predecessors 
    -- CP-element group 264: 	266 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	266 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u12_u12_553_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u12_u12_553_Update/cr
      -- CP-element group 264: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u12_u12_553_update_start_
      -- 
    -- logger for CP element group try1_CP_1680_elements(264)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(264)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(264) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_553_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(264), ack => ADD_u12_u12_553_inst_req_1); -- 
    try1_cp_element_group_264: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_264"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(144) & try1_CP_1680_elements(266);
      gj_try1_cp_element_group_264 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(264), clk => clk, reset => reset); --
    end block;
    -- CP-element group 265:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	263 
    -- CP-element group 265: successors 
    -- CP-element group 265: marked-successors 
    -- CP-element group 265: 	143 
    -- CP-element group 265: 	263 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u12_u12_553_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u12_u12_553_Sample/ra
      -- CP-element group 265: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u12_u12_553_sample_completed_
      -- 
    -- logger for CP element group try1_CP_1680_elements(265)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(265)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(265) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_553_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_553_inst_ack_0, ack => try1_CP_1680_elements(265)); -- 
    -- CP-element group 266:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	264 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	140 
    -- CP-element group 266: marked-successors 
    -- CP-element group 266: 	142 
    -- CP-element group 266: 	264 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u12_u12_553_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u12_u12_553_Update/ca
      -- CP-element group 266: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u12_u12_553_update_completed_
      -- 
    -- logger for CP element group try1_CP_1680_elements(266)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(266)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(266) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_553_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_553_inst_ack_1, ack => try1_CP_1680_elements(266)); -- 
    -- CP-element group 267:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	272 
    -- CP-element group 267: marked-predecessors 
    -- CP-element group 267: 	273 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	273 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_558_Sample/rr
      -- CP-element group 267: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_558_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_558_sample_start_
      -- 
    -- logger for CP element group try1_CP_1680_elements(267)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(267)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(267) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u16_u16_558_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(267), ack => ADD_u16_u16_558_inst_req_0); -- 
    try1_cp_element_group_267: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_267"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(272) & try1_CP_1680_elements(273);
      gj_try1_cp_element_group_267 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(267), clk => clk, reset => reset); --
    end block;
    -- CP-element group 268:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: marked-predecessors 
    -- CP-element group 268: 	274 
    -- CP-element group 268: 	277 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	274 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_558_update_start_
      -- CP-element group 268: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_558_Update/$entry
      -- CP-element group 268: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_558_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(268)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(268)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(268) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u16_u16_558_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(268), ack => ADD_u16_u16_558_inst_req_1); -- 
    try1_cp_element_group_268: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_268"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(274) & try1_CP_1680_elements(277);
      gj_try1_cp_element_group_268 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(268), clk => clk, reset => reset); --
    end block;
    -- CP-element group 269:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	139 
    -- CP-element group 269: marked-predecessors 
    -- CP-element group 269: 	271 
    -- CP-element group 269: 	277 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	271 
    -- CP-element group 269:  members (5) 
      -- CP-element group 269: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_Sample/word_access_start/$entry
      -- CP-element group 269: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_Sample/word_access_start/word_0/$entry
      -- CP-element group 269: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_Sample/word_access_start/word_0/rr
      -- CP-element group 269: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_sample_start_
      -- CP-element group 269: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_Sample/$entry
      -- 
    -- logger for CP element group try1_CP_1680_elements(269)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(269)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(269) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_PJ_556_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(269), ack => LOAD_PJ_556_load_0_req_0); -- 
    try1_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(139) & try1_CP_1680_elements(271) & try1_CP_1680_elements(277);
      gj_try1_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: marked-predecessors 
    -- CP-element group 270: 	272 
    -- CP-element group 270: 	273 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	272 
    -- CP-element group 270:  members (5) 
      -- CP-element group 270: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_update_start_
      -- CP-element group 270: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_Update/$entry
      -- CP-element group 270: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_Update/word_access_complete/word_0/cr
      -- CP-element group 270: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_Update/word_access_complete/word_0/$entry
      -- CP-element group 270: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_Update/word_access_complete/$entry
      -- 
    -- logger for CP element group try1_CP_1680_elements(270)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(270)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(270) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_PJ_556_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(270), ack => LOAD_PJ_556_load_0_req_1); -- 
    try1_cp_element_group_270: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_270"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(272) & try1_CP_1680_elements(273);
      gj_try1_cp_element_group_270 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(270), clk => clk, reset => reset); --
    end block;
    -- CP-element group 271:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	269 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	287 
    -- CP-element group 271: marked-successors 
    -- CP-element group 271: 	269 
    -- CP-element group 271:  members (5) 
      -- CP-element group 271: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_Sample/word_access_start/$exit
      -- CP-element group 271: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_Sample/word_access_start/word_0/$exit
      -- CP-element group 271: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_sample_completed_
      -- CP-element group 271: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_Sample/word_access_start/word_0/ra
      -- CP-element group 271: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_Sample/$exit
      -- 
    -- logger for CP element group try1_CP_1680_elements(271)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(271)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(271) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_PJ_556_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_PJ_556_load_0_ack_0, ack => try1_CP_1680_elements(271)); -- 
    -- CP-element group 272:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	270 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	267 
    -- CP-element group 272: marked-successors 
    -- CP-element group 272: 	270 
    -- CP-element group 272:  members (9) 
      -- CP-element group 272: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_Update/word_access_complete/word_0/ca
      -- CP-element group 272: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_Update/$exit
      -- CP-element group 272: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_Update/LOAD_PJ_556_Merge/merge_ack
      -- CP-element group 272: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_update_completed_
      -- CP-element group 272: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_Update/word_access_complete/word_0/$exit
      -- CP-element group 272: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_Update/LOAD_PJ_556_Merge/$entry
      -- CP-element group 272: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_Update/LOAD_PJ_556_Merge/$exit
      -- CP-element group 272: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_Update/LOAD_PJ_556_Merge/merge_req
      -- CP-element group 272: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_Update/word_access_complete/$exit
      -- 
    -- logger for CP element group try1_CP_1680_elements(272)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(272)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(272) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_PJ_556_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_PJ_556_load_0_ack_1, ack => try1_CP_1680_elements(272)); -- 
    -- CP-element group 273:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	267 
    -- CP-element group 273: successors 
    -- CP-element group 273: marked-successors 
    -- CP-element group 273: 	267 
    -- CP-element group 273: 	270 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_558_Sample/ra
      -- CP-element group 273: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_558_sample_completed_
      -- CP-element group 273: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_558_Sample/$exit
      -- 
    -- logger for CP element group try1_CP_1680_elements(273)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(273)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(273) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u16_u16_558_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_558_inst_ack_0, ack => try1_CP_1680_elements(273)); -- 
    -- CP-element group 274:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	268 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274: marked-successors 
    -- CP-element group 274: 	268 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_558_update_completed_
      -- CP-element group 274: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_558_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ADD_u16_u16_558_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(274)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(274)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(274) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u16_u16_558_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_558_inst_ack_1, ack => try1_CP_1680_elements(274)); -- 
    -- CP-element group 275:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	139 
    -- CP-element group 275: 	274 
    -- CP-element group 275: 	283 
    -- CP-element group 275: 	284 
    -- CP-element group 275: 	285 
    -- CP-element group 275: 	286 
    -- CP-element group 275: 	287 
    -- CP-element group 275: marked-predecessors 
    -- CP-element group 275: 	277 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	277 
    -- CP-element group 275:  members (9) 
      -- CP-element group 275: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_Sample/STORE_PJ_555_Split/$entry
      -- CP-element group 275: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_Sample/word_access_start/$entry
      -- CP-element group 275: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_Sample/STORE_PJ_555_Split/split_ack
      -- CP-element group 275: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_Sample/word_access_start/word_0/rr
      -- CP-element group 275: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_Sample/STORE_PJ_555_Split/$exit
      -- CP-element group 275: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_sample_start_
      -- CP-element group 275: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_Sample/STORE_PJ_555_Split/split_req
      -- CP-element group 275: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_Sample/$entry
      -- CP-element group 275: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_Sample/word_access_start/word_0/$entry
      -- 
    -- logger for CP element group try1_CP_1680_elements(275)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(275)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(275) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:STORE_PJ_555_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(275), ack => STORE_PJ_555_store_0_req_0); -- 
    try1_cp_element_group_275: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_275"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= try1_CP_1680_elements(139) & try1_CP_1680_elements(274) & try1_CP_1680_elements(283) & try1_CP_1680_elements(284) & try1_CP_1680_elements(285) & try1_CP_1680_elements(286) & try1_CP_1680_elements(287) & try1_CP_1680_elements(277);
      gj_try1_cp_element_group_275 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(275), clk => clk, reset => reset); --
    end block;
    -- CP-element group 276:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: marked-predecessors 
    -- CP-element group 276: 	278 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	278 
    -- CP-element group 276:  members (5) 
      -- CP-element group 276: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_Update/word_access_complete/$entry
      -- CP-element group 276: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_Update/word_access_complete/word_0/$entry
      -- CP-element group 276: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_Update/word_access_complete/word_0/cr
      -- CP-element group 276: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_update_start_
      -- CP-element group 276: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_Update/$entry
      -- 
    -- logger for CP element group try1_CP_1680_elements(276)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(276)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(276) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:STORE_PJ_555_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(276), ack => STORE_PJ_555_store_0_req_1); -- 
    try1_cp_element_group_276: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_276"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(278);
      gj_try1_cp_element_group_276 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(276), clk => clk, reset => reset); --
    end block;
    -- CP-element group 277:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	275 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	288 
    -- CP-element group 277: marked-successors 
    -- CP-element group 277: 	201 
    -- CP-element group 277: 	268 
    -- CP-element group 277: 	269 
    -- CP-element group 277: 	275 
    -- CP-element group 277: 	207 
    -- CP-element group 277: 	233 
    -- CP-element group 277: 	241 
    -- CP-element group 277:  members (6) 
      -- CP-element group 277: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_Sample/word_access_start/$exit
      -- CP-element group 277: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_Sample/word_access_start/word_0/ra
      -- CP-element group 277: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_sample_completed_
      -- CP-element group 277: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_Sample/word_access_start/word_0/$exit
      -- CP-element group 277: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/ring_reenable_memory_space_0
      -- 
    -- logger for CP element group try1_CP_1680_elements(277)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(277)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(277) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:STORE_PJ_555_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_PJ_555_store_0_ack_0, ack => try1_CP_1680_elements(277)); -- 
    -- CP-element group 278:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	276 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	288 
    -- CP-element group 278: marked-successors 
    -- CP-element group 278: 	276 
    -- CP-element group 278:  members (5) 
      -- CP-element group 278: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_Update/word_access_complete/$exit
      -- CP-element group 278: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_Update/word_access_complete/word_0/$exit
      -- CP-element group 278: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_update_completed_
      -- CP-element group 278: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/STORE_PJ_555_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(278)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(278)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(278) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:STORE_PJ_555_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_PJ_555_store_0_ack_1, ack => try1_CP_1680_elements(278)); -- 
    -- CP-element group 279:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	139 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	140 
    -- CP-element group 279:  members (1) 
      -- CP-element group 279: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group try1_CP_1680_elements(279)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(279)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(279) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(279) is a control-delay.
    cp_element_279_delay: control_delay_element  generic map(name => " 279_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(139), ack => try1_CP_1680_elements(279), clk => clk, reset =>reset);
    -- CP-element group 280:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	213 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	219 
    -- CP-element group 280:  members (1) 
      -- CP-element group 280: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_508_array_obj_ref_515_delay
      -- 
    -- logger for CP element group try1_CP_1680_elements(280)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(280)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(280) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(280) is a control-delay.
    cp_element_280_delay: control_delay_element  generic map(name => " 280_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(213), ack => try1_CP_1680_elements(280), clk => clk, reset =>reset);
    -- CP-element group 281:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	221 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	251 
    -- CP-element group 281:  members (1) 
      -- CP-element group 281: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_515_array_obj_ref_540_delay
      -- 
    -- logger for CP element group try1_CP_1680_elements(281)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(281)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(281) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(281) is a control-delay.
    cp_element_281_delay: control_delay_element  generic map(name => " 281_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(221), ack => try1_CP_1680_elements(281), clk => clk, reset =>reset);
    -- CP-element group 282:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	253 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	259 
    -- CP-element group 282:  members (1) 
      -- CP-element group 282: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/array_obj_ref_540_array_obj_ref_547_delay
      -- 
    -- logger for CP element group try1_CP_1680_elements(282)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(282)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(282) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(282) is a control-delay.
    cp_element_282_delay: control_delay_element  generic map(name => " 282_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(253), ack => try1_CP_1680_elements(282), clk => clk, reset =>reset);
    -- CP-element group 283:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	203 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	275 
    -- CP-element group 283:  members (1) 
      -- CP-element group 283: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_500_STORE_PJ_555_delay
      -- 
    -- logger for CP element group try1_CP_1680_elements(283)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(283)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(283) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(283) is a control-delay.
    cp_element_283_delay: control_delay_element  generic map(name => " 283_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(203), ack => try1_CP_1680_elements(283), clk => clk, reset =>reset);
    -- CP-element group 284:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	209 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	275 
    -- CP-element group 284:  members (1) 
      -- CP-element group 284: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_505_STORE_PJ_555_delay
      -- 
    -- logger for CP element group try1_CP_1680_elements(284)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(284)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(284) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(284) is a control-delay.
    cp_element_284_delay: control_delay_element  generic map(name => " 284_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(209), ack => try1_CP_1680_elements(284), clk => clk, reset =>reset);
    -- CP-element group 285:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	235 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	275 
    -- CP-element group 285:  members (1) 
      -- CP-element group 285: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_527_STORE_PJ_555_delay
      -- 
    -- logger for CP element group try1_CP_1680_elements(285)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(285)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(285) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(285) is a control-delay.
    cp_element_285_delay: control_delay_element  generic map(name => " 285_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(235), ack => try1_CP_1680_elements(285), clk => clk, reset =>reset);
    -- CP-element group 286:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	243 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	275 
    -- CP-element group 286:  members (1) 
      -- CP-element group 286: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_532_STORE_PJ_555_delay
      -- 
    -- logger for CP element group try1_CP_1680_elements(286)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(286)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(286) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(286) is a control-delay.
    cp_element_286_delay: control_delay_element  generic map(name => " 286_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(243), ack => try1_CP_1680_elements(286), clk => clk, reset =>reset);
    -- CP-element group 287:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	271 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	275 
    -- CP-element group 287:  members (1) 
      -- CP-element group 287: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/LOAD_PJ_556_STORE_PJ_555_delay
      -- 
    -- logger for CP element group try1_CP_1680_elements(287)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(287)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(287) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(287) is a control-delay.
    cp_element_287_delay: control_delay_element  generic map(name => " 287_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(271), ack => try1_CP_1680_elements(287), clk => clk, reset =>reset);
    -- CP-element group 288:  join  transition  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	254 
    -- CP-element group 288: 	261 
    -- CP-element group 288: 	262 
    -- CP-element group 288: 	277 
    -- CP-element group 288: 	214 
    -- CP-element group 288: 	278 
    -- CP-element group 288: 	222 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	136 
    -- CP-element group 288:  members (1) 
      -- CP-element group 288: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/do_while_stmt_455_loop_body/$exit
      -- 
    -- logger for CP element group try1_CP_1680_elements(288)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(288)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(288) fired."); 
        -- 
      end if; --
    end process; 
    try1_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= try1_CP_1680_elements(254) & try1_CP_1680_elements(261) & try1_CP_1680_elements(262) & try1_CP_1680_elements(277) & try1_CP_1680_elements(214) & try1_CP_1680_elements(278) & try1_CP_1680_elements(222);
      gj_try1_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  transition  input  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	135 
    -- CP-element group 289: successors 
    -- CP-element group 289:  members (2) 
      -- CP-element group 289: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/loop_exit/$exit
      -- CP-element group 289: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/loop_exit/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(289)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(289)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(289) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:do_while_stmt_455_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_455_branch_ack_0, ack => try1_CP_1680_elements(289)); -- 
    -- CP-element group 290:  transition  input  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	135 
    -- CP-element group 290: successors 
    -- CP-element group 290:  members (2) 
      -- CP-element group 290: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/loop_taken/$exit
      -- CP-element group 290: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/loop_taken/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(290)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(290)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(290) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:do_while_stmt_455_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_455_branch_ack_1, ack => try1_CP_1680_elements(290)); -- 
    -- CP-element group 291:  transition  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	133 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	131 
    -- CP-element group 291:  members (1) 
      -- CP-element group 291: 	 branch_block_stmt_443/branch_block_stmt_454/do_while_stmt_455/$exit
      -- 
    -- logger for CP element group try1_CP_1680_elements(291)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(291)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(291) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(291) <= try1_CP_1680_elements(133);
    -- CP-element group 292:  transition  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	517 
    -- CP-element group 292: successors 
    -- CP-element group 292:  members (5) 
      -- CP-element group 292: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_sample_completed_
      -- CP-element group 292: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_Sample/$exit
      -- CP-element group 292: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_Sample/word_access_start/$exit
      -- CP-element group 292: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_Sample/word_access_start/word_0/$exit
      -- CP-element group 292: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(292)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(292)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(292) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:STORE_total_573_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_total_573_store_0_ack_0, ack => try1_CP_1680_elements(292)); -- 
    -- CP-element group 293:  transition  place  input  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	517 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	295 
    -- CP-element group 293:  members (11) 
      -- CP-element group 293: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575__exit__
      -- CP-element group 293: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576__entry__
      -- CP-element group 293: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/branch_block_stmt_576__entry__
      -- CP-element group 293: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577__entry__
      -- CP-element group 293: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/$exit
      -- CP-element group 293: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_update_completed_
      -- CP-element group 293: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_Update/$exit
      -- CP-element group 293: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_Update/word_access_complete/$exit
      -- CP-element group 293: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_Update/word_access_complete/word_0/$exit
      -- CP-element group 293: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_Update/word_access_complete/word_0/ca
      -- CP-element group 293: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/$entry
      -- 
    -- logger for CP element group try1_CP_1680_elements(293)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(293)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(293) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:STORE_total_573_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_total_573_store_0_ack_1, ack => try1_CP_1680_elements(293)); -- 
    -- CP-element group 294:  fork  transition  place  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	369 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	385 
    -- CP-element group 294: 	377 
    -- CP-element group 294: 	378 
    -- CP-element group 294: 	380 
    -- CP-element group 294: 	371 
    -- CP-element group 294: 	372 
    -- CP-element group 294: 	373 
    -- CP-element group 294: 	374 
    -- CP-element group 294: 	376 
    -- CP-element group 294:  members (47) 
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577__exit__
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576__exit__
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638__entry__
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/branch_block_stmt_576__exit__
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/$exit
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/$entry
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/call_stmt_624_update_start_
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/ADD_u12_u12_621_sample_start_
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/ADD_u12_u12_621_update_start_
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/ADD_u12_u12_621_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/ADD_u12_u12_621_Sample/rr
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/ADD_u12_u12_621_Update/$entry
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/ADD_u12_u12_621_Update/cr
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_sample_start_
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_update_start_
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_word_address_calculated
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_root_address_calculated
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_Sample/word_access_start/$entry
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_Sample/word_access_start/word_0/$entry
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_Sample/word_access_start/word_0/rr
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_Update/$entry
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_Update/word_access_complete/$entry
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_Update/word_access_complete/word_0/$entry
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_Update/word_access_complete/word_0/cr
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/call_stmt_624_Update/$entry
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/call_stmt_624_Update/ccr
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/CONCAT_u4_u16_630_update_start_
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_sample_start_
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_update_start_
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_word_address_calculated
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_root_address_calculated
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_Sample/word_access_start/$entry
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_Sample/word_access_start/word_0/$entry
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_Sample/word_access_start/word_0/rr
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_Update/$entry
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_Update/word_access_complete/$entry
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_Update/word_access_complete/word_0/$entry
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_Update/word_access_complete/word_0/cr
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/CONCAT_u4_u16_630_Update/$entry
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/CONCAT_u4_u16_630_Update/cr
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_update_start_
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_Update/$entry
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_Update/word_access_complete/$entry
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_Update/word_access_complete/word_0/$entry
      -- CP-element group 294: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(294)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(294)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(294) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_621_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_621_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_total_622_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_total_622_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:call_stmt_624_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_zer_626_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_zer_626_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:CONCAT_u4_u16_630_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_637_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    rr_3736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(294), ack => ADD_u12_u12_621_inst_req_0); -- 
    cr_3741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(294), ack => ADD_u12_u12_621_inst_req_1); -- 
    rr_3758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(294), ack => LOAD_total_622_load_0_req_0); -- 
    cr_3769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(294), ack => LOAD_total_622_load_0_req_1); -- 
    ccr_3784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(294), ack => call_stmt_624_call_req_1); -- 
    rr_3805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(294), ack => LOAD_zer_626_load_0_req_0); -- 
    cr_3816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(294), ack => LOAD_zer_626_load_0_req_1); -- 
    cr_3831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(294), ack => CONCAT_u4_u16_630_inst_req_1); -- 
    cr_3903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(294), ack => array_obj_ref_637_load_0_req_1); -- 
    try1_CP_1680_elements(294) <= try1_CP_1680_elements(369);
    -- CP-element group 295:  transition  place  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	293 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	301 
    -- CP-element group 295:  members (2) 
      -- CP-element group 295: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577__entry__
      -- CP-element group 295: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/$entry
      -- 
    -- logger for CP element group try1_CP_1680_elements(295)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(295)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(295) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(295) <= try1_CP_1680_elements(293);
    -- CP-element group 296:  merge  place  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	369 
    -- CP-element group 296:  members (1) 
      -- CP-element group 296: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577__exit__
      -- 
    -- logger for CP element group try1_CP_1680_elements(296)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(296)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(296) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(296) is bound as output of CP function.
    -- CP-element group 297:  merge  place  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	300 
    -- CP-element group 297:  members (1) 
      -- CP-element group 297: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/loop_back
      -- 
    -- logger for CP element group try1_CP_1680_elements(297)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(297)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(297) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(297) is bound as output of CP function.
    -- CP-element group 298:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	303 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	367 
    -- CP-element group 298: 	368 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/condition_done
      -- CP-element group 298: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/loop_exit/$entry
      -- CP-element group 298: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/loop_taken/$entry
      -- 
    -- logger for CP element group try1_CP_1680_elements(298)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(298)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(298) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(298) <= try1_CP_1680_elements(303);
    -- CP-element group 299:  branch  place  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	366 
    -- CP-element group 299: successors 
    -- CP-element group 299:  members (1) 
      -- CP-element group 299: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/loop_body_done
      -- 
    -- logger for CP element group try1_CP_1680_elements(299)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(299)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(299) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(299) <= try1_CP_1680_elements(366);
    -- CP-element group 300:  transition  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	297 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	309 
    -- CP-element group 300:  members (1) 
      -- CP-element group 300: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group try1_CP_1680_elements(300)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(300)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(300) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(300) <= try1_CP_1680_elements(297);
    -- CP-element group 301:  transition  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	295 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	311 
    -- CP-element group 301:  members (1) 
      -- CP-element group 301: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group try1_CP_1680_elements(301)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(301)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(301) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(301) <= try1_CP_1680_elements(295);
    -- CP-element group 302:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	305 
    -- CP-element group 302: 	306 
    -- CP-element group 302: 	344 
    -- CP-element group 302: 	354 
    -- CP-element group 302: 	362 
    -- CP-element group 302:  members (6) 
      -- CP-element group 302: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/$entry
      -- CP-element group 302: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/loop_body_start
      -- CP-element group 302: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_word_address_calculated
      -- CP-element group 302: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_root_address_calculated
      -- CP-element group 302: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_word_address_calculated
      -- CP-element group 302: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_root_address_calculated
      -- 
    -- logger for CP element group try1_CP_1680_elements(302)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(302)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(302) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(302) is bound as output of CP function.
    -- CP-element group 303:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	308 
    -- CP-element group 303: 	361 
    -- CP-element group 303: 	362 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	298 
    -- CP-element group 303:  members (1) 
      -- CP-element group 303: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/condition_evaluated
      -- 
    -- logger for CP element group try1_CP_1680_elements(303)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(303)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(303) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:do_while_stmt_577_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_3285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(303), ack => do_while_stmt_577_branch_req_0); -- 
    try1_cp_element_group_303: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_303"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(308) & try1_CP_1680_elements(361) & try1_CP_1680_elements(362);
      gj_try1_cp_element_group_303 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(303), clk => clk, reset => reset); --
    end block;
    -- CP-element group 304:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	305 
    -- CP-element group 304: marked-predecessors 
    -- CP-element group 304: 	308 
    -- CP-element group 304: successors 
    -- CP-element group 304:  members (2) 
      -- CP-element group 304: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/aggregated_phi_sample_req
      -- CP-element group 304: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/phi_stmt_579_sample_start__ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(304)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(304)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(304) fired."); 
        -- 
      end if; --
    end process; 
    try1_cp_element_group_304: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_304"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(305) & try1_CP_1680_elements(308);
      gj_try1_cp_element_group_304 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(304), clk => clk, reset => reset); --
    end block;
    -- CP-element group 305:  join  transition  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	302 
    -- CP-element group 305: marked-predecessors 
    -- CP-element group 305: 	307 
    -- CP-element group 305: 	361 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	304 
    -- CP-element group 305:  members (1) 
      -- CP-element group 305: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/phi_stmt_579_sample_start_
      -- 
    -- logger for CP element group try1_CP_1680_elements(305)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(305)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(305) fired."); 
        -- 
      end if; --
    end process; 
    try1_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(302) & try1_CP_1680_elements(307) & try1_CP_1680_elements(361);
      gj_try1_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	302 
    -- CP-element group 306: marked-predecessors 
    -- CP-element group 306: 	308 
    -- CP-element group 306: 	324 
    -- CP-element group 306: 	328 
    -- CP-element group 306: 	332 
    -- CP-element group 306: 	350 
    -- CP-element group 306: 	360 
    -- CP-element group 306: successors 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/aggregated_phi_update_req
      -- CP-element group 306: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/phi_stmt_579_update_start_
      -- CP-element group 306: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/phi_stmt_579_update_start__ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(306)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(306)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(306) fired."); 
        -- 
      end if; --
    end process; 
    try1_cp_element_group_306: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_306"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= try1_CP_1680_elements(302) & try1_CP_1680_elements(308) & try1_CP_1680_elements(324) & try1_CP_1680_elements(328) & try1_CP_1680_elements(332) & try1_CP_1680_elements(350) & try1_CP_1680_elements(360);
      gj_try1_cp_element_group_306 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(306), clk => clk, reset => reset); --
    end block;
    -- CP-element group 307:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	359 
    -- CP-element group 307: marked-successors 
    -- CP-element group 307: 	305 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/aggregated_phi_sample_ack
      -- CP-element group 307: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/phi_stmt_579_sample_completed_
      -- CP-element group 307: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/phi_stmt_579_sample_completed__ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(307)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(307)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(307) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(307) is bound as output of CP function.
    -- CP-element group 308:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	303 
    -- CP-element group 308: 	322 
    -- CP-element group 308: 	326 
    -- CP-element group 308: 	330 
    -- CP-element group 308: 	348 
    -- CP-element group 308: 	358 
    -- CP-element group 308: marked-successors 
    -- CP-element group 308: 	304 
    -- CP-element group 308: 	306 
    -- CP-element group 308:  members (81) 
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/aggregated_phi_update_ack
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/phi_stmt_579_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/phi_stmt_579_update_completed__ps
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_word_address_calculated
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_root_address_calculated
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_offset_calculated
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_index_resized_0
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_index_scaled_0
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_index_computed_0
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_index_resize_0/$entry
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_index_resize_0/$exit
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_index_resize_0/index_resize_req
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_index_resize_0/index_resize_ack
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_index_scale_0/$entry
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_index_scale_0/$exit
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_index_scale_0/scale_rename_req
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_index_scale_0/scale_rename_ack
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_final_index_sum_regn/$entry
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_final_index_sum_regn/$exit
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_final_index_sum_regn/req
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_final_index_sum_regn/ack
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_base_plus_offset/$entry
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_base_plus_offset/$exit
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_base_plus_offset/sum_rename_req
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_base_plus_offset/sum_rename_ack
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_word_addrgen/$entry
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_word_addrgen/$exit
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_word_addrgen/root_register_req
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_word_addrgen/root_register_ack
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_index_scaled_0
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_word_address_calculated
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_root_address_calculated
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_offset_calculated
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_index_resized_0
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_index_scaled_0
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_index_computed_0
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_index_resize_0/$entry
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_index_resize_0/$exit
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_index_resize_0/index_resize_req
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_index_resize_0/index_resize_ack
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_index_scale_0/$entry
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_index_scale_0/$exit
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_index_scale_0/scale_rename_req
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_index_scale_0/scale_rename_ack
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_final_index_sum_regn/$entry
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_final_index_sum_regn/$exit
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_final_index_sum_regn/req
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_final_index_sum_regn/ack
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_base_plus_offset/$entry
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_base_plus_offset/$exit
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_base_plus_offset/sum_rename_req
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_base_plus_offset/sum_rename_ack
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_word_addrgen/$entry
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_word_addrgen/$exit
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_word_addrgen/root_register_req
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_word_addrgen/root_register_ack
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_word_address_calculated
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_root_address_calculated
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_offset_calculated
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_index_resized_0
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_index_computed_0
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_index_resize_0/$entry
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_index_resize_0/$exit
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_index_resize_0/index_resize_req
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_index_resize_0/index_resize_ack
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_index_scale_0/$entry
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_index_scale_0/$exit
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_index_scale_0/scale_rename_req
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_index_scale_0/scale_rename_ack
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_final_index_sum_regn/$entry
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_final_index_sum_regn/$exit
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_final_index_sum_regn/req
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_final_index_sum_regn/ack
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_base_plus_offset/$entry
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_base_plus_offset/$exit
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_base_plus_offset/sum_rename_req
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_base_plus_offset/sum_rename_ack
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_word_addrgen/$entry
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_word_addrgen/$exit
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_word_addrgen/root_register_req
      -- CP-element group 308: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(308)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(308)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(308) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(308) is bound as output of CP function.
    -- CP-element group 309:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	300 
    -- CP-element group 309: successors 
    -- CP-element group 309:  members (1) 
      -- CP-element group 309: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/phi_stmt_579_loopback_trigger
      -- 
    -- logger for CP element group try1_CP_1680_elements(309)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(309)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(309) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(309) <= try1_CP_1680_elements(300);
    -- CP-element group 310:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: successors 
    -- CP-element group 310:  members (2) 
      -- CP-element group 310: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/phi_stmt_579_loopback_sample_req
      -- CP-element group 310: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/phi_stmt_579_loopback_sample_req_ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(310)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(310)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(310) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:phi_stmt_579_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_579_loopback_sample_req_3300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_579_loopback_sample_req_3300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(310), ack => phi_stmt_579_req_1); -- 
    -- Element group try1_CP_1680_elements(310) is bound as output of CP function.
    -- CP-element group 311:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	301 
    -- CP-element group 311: successors 
    -- CP-element group 311:  members (1) 
      -- CP-element group 311: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/phi_stmt_579_entry_trigger
      -- 
    -- logger for CP element group try1_CP_1680_elements(311)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(311)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(311) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(311) <= try1_CP_1680_elements(301);
    -- CP-element group 312:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: successors 
    -- CP-element group 312:  members (2) 
      -- CP-element group 312: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/phi_stmt_579_entry_sample_req
      -- CP-element group 312: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/phi_stmt_579_entry_sample_req_ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(312)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(312)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(312) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:phi_stmt_579_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_579_entry_sample_req_3303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_579_entry_sample_req_3303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(312), ack => phi_stmt_579_req_0); -- 
    -- Element group try1_CP_1680_elements(312) is bound as output of CP function.
    -- CP-element group 313:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: successors 
    -- CP-element group 313:  members (2) 
      -- CP-element group 313: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/phi_stmt_579_phi_mux_ack
      -- CP-element group 313: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/phi_stmt_579_phi_mux_ack_ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(313)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(313)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(313) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:phi_stmt_579_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_579_phi_mux_ack_3306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_579_ack_0, ack => try1_CP_1680_elements(313)); -- 
    -- CP-element group 314:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: successors 
    -- CP-element group 314:  members (4) 
      -- CP-element group 314: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/type_cast_582_sample_start__ps
      -- CP-element group 314: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/type_cast_582_sample_completed__ps
      -- CP-element group 314: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/type_cast_582_sample_start_
      -- CP-element group 314: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/type_cast_582_sample_completed_
      -- 
    -- logger for CP element group try1_CP_1680_elements(314)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(314)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(314) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(314) is bound as output of CP function.
    -- CP-element group 315:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	317 
    -- CP-element group 315:  members (2) 
      -- CP-element group 315: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/type_cast_582_update_start__ps
      -- CP-element group 315: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/type_cast_582_update_start_
      -- 
    -- logger for CP element group try1_CP_1680_elements(315)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(315)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(315) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(315) is bound as output of CP function.
    -- CP-element group 316:  join  transition  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	317 
    -- CP-element group 316: successors 
    -- CP-element group 316:  members (1) 
      -- CP-element group 316: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/type_cast_582_update_completed__ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(316)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(316)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(316) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(316) <= try1_CP_1680_elements(317);
    -- CP-element group 317:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	315 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	316 
    -- CP-element group 317:  members (1) 
      -- CP-element group 317: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/type_cast_582_update_completed_
      -- 
    -- logger for CP element group try1_CP_1680_elements(317)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(317)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(317) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(317) is a control-delay.
    cp_element_317_delay: control_delay_element  generic map(name => " 317_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(315), ack => try1_CP_1680_elements(317), clk => clk, reset =>reset);
    -- CP-element group 318:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	320 
    -- CP-element group 318:  members (4) 
      -- CP-element group 318: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/R_NK_583_sample_start__ps
      -- CP-element group 318: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/R_NK_583_sample_start_
      -- CP-element group 318: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/R_NK_583_Sample/$entry
      -- CP-element group 318: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/R_NK_583_Sample/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(318)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(318)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(318) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NK_612_583_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(318), ack => NK_612_583_buf_req_0); -- 
    -- Element group try1_CP_1680_elements(318) is bound as output of CP function.
    -- CP-element group 319:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	321 
    -- CP-element group 319:  members (4) 
      -- CP-element group 319: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/R_NK_583_update_start__ps
      -- CP-element group 319: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/R_NK_583_update_start_
      -- CP-element group 319: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/R_NK_583_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/R_NK_583_Update/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(319)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(319)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(319) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NK_612_583_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(319), ack => NK_612_583_buf_req_1); -- 
    -- Element group try1_CP_1680_elements(319) is bound as output of CP function.
    -- CP-element group 320:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	318 
    -- CP-element group 320: successors 
    -- CP-element group 320:  members (4) 
      -- CP-element group 320: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/R_NK_583_sample_completed__ps
      -- CP-element group 320: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/R_NK_583_sample_completed_
      -- CP-element group 320: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/R_NK_583_Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/R_NK_583_Sample/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(320)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(320)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(320) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NK_612_583_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NK_612_583_buf_ack_0, ack => try1_CP_1680_elements(320)); -- 
    -- CP-element group 321:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	319 
    -- CP-element group 321: successors 
    -- CP-element group 321:  members (4) 
      -- CP-element group 321: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/R_NK_583_update_completed__ps
      -- CP-element group 321: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/R_NK_583_update_completed_
      -- CP-element group 321: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/R_NK_583_Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/R_NK_583_Update/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(321)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(321)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(321) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NK_612_583_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NK_612_583_buf_ack_1, ack => try1_CP_1680_elements(321)); -- 
    -- CP-element group 322:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	308 
    -- CP-element group 322: marked-predecessors 
    -- CP-element group 322: 	324 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	324 
    -- CP-element group 322:  members (5) 
      -- CP-element group 322: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_sample_start_
      -- CP-element group 322: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_Sample/word_access_start/$entry
      -- CP-element group 322: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_Sample/word_access_start/word_0/$entry
      -- CP-element group 322: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(322)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(322)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(322) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_587_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(322), ack => array_obj_ref_587_load_0_req_0); -- 
    try1_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(308) & try1_CP_1680_elements(324);
      gj_try1_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: marked-predecessors 
    -- CP-element group 323: 	325 
    -- CP-element group 323: 	336 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	325 
    -- CP-element group 323:  members (5) 
      -- CP-element group 323: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_update_start_
      -- CP-element group 323: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_Update/word_access_complete/$entry
      -- CP-element group 323: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_Update/word_access_complete/word_0/$entry
      -- CP-element group 323: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(323)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(323)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(323) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_587_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(323), ack => array_obj_ref_587_load_0_req_1); -- 
    try1_cp_element_group_323: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_323"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(325) & try1_CP_1680_elements(336);
      gj_try1_cp_element_group_323 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(323), clk => clk, reset => reset); --
    end block;
    -- CP-element group 324:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	322 
    -- CP-element group 324: successors 
    -- CP-element group 324: marked-successors 
    -- CP-element group 324: 	306 
    -- CP-element group 324: 	322 
    -- CP-element group 324:  members (5) 
      -- CP-element group 324: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_sample_completed_
      -- CP-element group 324: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_Sample/$exit
      -- CP-element group 324: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_Sample/word_access_start/$exit
      -- CP-element group 324: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_Sample/word_access_start/word_0/$exit
      -- CP-element group 324: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(324)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(324)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(324) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_587_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_587_load_0_ack_0, ack => try1_CP_1680_elements(324)); -- 
    -- CP-element group 325:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	323 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	334 
    -- CP-element group 325: marked-successors 
    -- CP-element group 325: 	323 
    -- CP-element group 325:  members (9) 
      -- CP-element group 325: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_update_completed_
      -- CP-element group 325: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_Update/$exit
      -- CP-element group 325: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_Update/word_access_complete/$exit
      -- CP-element group 325: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_Update/word_access_complete/word_0/$exit
      -- CP-element group 325: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_Update/word_access_complete/word_0/ca
      -- CP-element group 325: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_Update/array_obj_ref_587_Merge/$entry
      -- CP-element group 325: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_Update/array_obj_ref_587_Merge/$exit
      -- CP-element group 325: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_Update/array_obj_ref_587_Merge/merge_req
      -- CP-element group 325: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_587_Update/array_obj_ref_587_Merge/merge_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(325)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(325)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(325) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_587_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_587_load_0_ack_1, ack => try1_CP_1680_elements(325)); -- 
    -- CP-element group 326:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	308 
    -- CP-element group 326: marked-predecessors 
    -- CP-element group 326: 	328 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	328 
    -- CP-element group 326:  members (5) 
      -- CP-element group 326: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_Sample/word_access_start/$entry
      -- CP-element group 326: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_Sample/word_access_start/word_0/$entry
      -- CP-element group 326: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(326)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(326)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(326) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_591_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(326), ack => array_obj_ref_591_load_0_req_0); -- 
    try1_cp_element_group_326: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_326"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(308) & try1_CP_1680_elements(328);
      gj_try1_cp_element_group_326 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(326), clk => clk, reset => reset); --
    end block;
    -- CP-element group 327:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: marked-predecessors 
    -- CP-element group 327: 	329 
    -- CP-element group 327: 	336 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	329 
    -- CP-element group 327:  members (5) 
      -- CP-element group 327: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_update_start_
      -- CP-element group 327: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_Update/$entry
      -- CP-element group 327: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_Update/word_access_complete/$entry
      -- CP-element group 327: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_Update/word_access_complete/word_0/$entry
      -- CP-element group 327: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(327)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(327)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(327) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_591_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(327), ack => array_obj_ref_591_load_0_req_1); -- 
    try1_cp_element_group_327: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_327"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(329) & try1_CP_1680_elements(336);
      gj_try1_cp_element_group_327 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(327), clk => clk, reset => reset); --
    end block;
    -- CP-element group 328:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	326 
    -- CP-element group 328: successors 
    -- CP-element group 328: marked-successors 
    -- CP-element group 328: 	306 
    -- CP-element group 328: 	326 
    -- CP-element group 328:  members (5) 
      -- CP-element group 328: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_sample_completed_
      -- CP-element group 328: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_Sample/$exit
      -- CP-element group 328: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_Sample/word_access_start/$exit
      -- CP-element group 328: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_Sample/word_access_start/word_0/$exit
      -- CP-element group 328: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(328)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(328)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(328) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_591_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_591_load_0_ack_0, ack => try1_CP_1680_elements(328)); -- 
    -- CP-element group 329:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	327 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	334 
    -- CP-element group 329: marked-successors 
    -- CP-element group 329: 	327 
    -- CP-element group 329:  members (9) 
      -- CP-element group 329: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_update_completed_
      -- CP-element group 329: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_Update/$exit
      -- CP-element group 329: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_Update/word_access_complete/$exit
      -- CP-element group 329: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_Update/word_access_complete/word_0/$exit
      -- CP-element group 329: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_Update/word_access_complete/word_0/ca
      -- CP-element group 329: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_Update/array_obj_ref_591_Merge/$entry
      -- CP-element group 329: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_Update/array_obj_ref_591_Merge/$exit
      -- CP-element group 329: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_Update/array_obj_ref_591_Merge/merge_req
      -- CP-element group 329: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_591_Update/array_obj_ref_591_Merge/merge_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(329)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(329)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(329) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_591_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_591_load_0_ack_1, ack => try1_CP_1680_elements(329)); -- 
    -- CP-element group 330:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	308 
    -- CP-element group 330: marked-predecessors 
    -- CP-element group 330: 	332 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	332 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/assign_stmt_595_sample_start_
      -- CP-element group 330: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/assign_stmt_595_Sample/$entry
      -- CP-element group 330: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/assign_stmt_595_Sample/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(330)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(330)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(330) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_K_517_delayed_5_0_593_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(330), ack => W_K_517_delayed_5_0_593_inst_req_0); -- 
    try1_cp_element_group_330: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_330"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(308) & try1_CP_1680_elements(332);
      gj_try1_cp_element_group_330 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(330), clk => clk, reset => reset); --
    end block;
    -- CP-element group 331:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: marked-predecessors 
    -- CP-element group 331: 	333 
    -- CP-element group 331: 	340 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	333 
    -- CP-element group 331:  members (3) 
      -- CP-element group 331: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/assign_stmt_595_update_start_
      -- CP-element group 331: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/assign_stmt_595_Update/$entry
      -- CP-element group 331: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/assign_stmt_595_Update/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(331)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(331)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(331) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_K_517_delayed_5_0_593_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(331), ack => W_K_517_delayed_5_0_593_inst_req_1); -- 
    try1_cp_element_group_331: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_331"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(333) & try1_CP_1680_elements(340);
      gj_try1_cp_element_group_331 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(331), clk => clk, reset => reset); --
    end block;
    -- CP-element group 332:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	330 
    -- CP-element group 332: successors 
    -- CP-element group 332: marked-successors 
    -- CP-element group 332: 	306 
    -- CP-element group 332: 	330 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/assign_stmt_595_sample_completed_
      -- CP-element group 332: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/assign_stmt_595_Sample/$exit
      -- CP-element group 332: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/assign_stmt_595_Sample/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(332)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(332)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(332) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_K_517_delayed_5_0_593_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K_517_delayed_5_0_593_inst_ack_0, ack => try1_CP_1680_elements(332)); -- 
    -- CP-element group 333:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	331 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	338 
    -- CP-element group 333: marked-successors 
    -- CP-element group 333: 	331 
    -- CP-element group 333:  members (29) 
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/assign_stmt_595_update_completed_
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/assign_stmt_595_Update/$exit
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/assign_stmt_595_Update/ack
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_word_address_calculated
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_root_address_calculated
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_offset_calculated
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_index_resized_0
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_index_scaled_0
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_index_computed_0
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_index_resize_0/$entry
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_index_resize_0/$exit
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_index_resize_0/index_resize_req
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_index_resize_0/index_resize_ack
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_index_scale_0/$entry
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_index_scale_0/$exit
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_index_scale_0/scale_rename_req
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_index_scale_0/scale_rename_ack
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_final_index_sum_regn/$entry
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_final_index_sum_regn/$exit
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_final_index_sum_regn/req
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_final_index_sum_regn/ack
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_base_plus_offset/$entry
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_base_plus_offset/$exit
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_base_plus_offset/sum_rename_req
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_base_plus_offset/sum_rename_ack
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_word_addrgen/$entry
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_word_addrgen/$exit
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_word_addrgen/root_register_req
      -- CP-element group 333: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(333)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(333)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(333) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_K_517_delayed_5_0_593_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_K_517_delayed_5_0_593_inst_ack_1, ack => try1_CP_1680_elements(333)); -- 
    -- CP-element group 334:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	325 
    -- CP-element group 334: 	329 
    -- CP-element group 334: marked-predecessors 
    -- CP-element group 334: 	336 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	336 
    -- CP-element group 334:  members (3) 
      -- CP-element group 334: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/MUL_u16_u16_600_sample_start_
      -- CP-element group 334: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/MUL_u16_u16_600_Sample/$entry
      -- CP-element group 334: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/MUL_u16_u16_600_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(334)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(334)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(334) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:MUL_u16_u16_600_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(334), ack => MUL_u16_u16_600_inst_req_0); -- 
    try1_cp_element_group_334: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_334"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(325) & try1_CP_1680_elements(329) & try1_CP_1680_elements(336);
      gj_try1_cp_element_group_334 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(334), clk => clk, reset => reset); --
    end block;
    -- CP-element group 335:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: marked-predecessors 
    -- CP-element group 335: 	337 
    -- CP-element group 335: 	340 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	337 
    -- CP-element group 335:  members (3) 
      -- CP-element group 335: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/MUL_u16_u16_600_update_start_
      -- CP-element group 335: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/MUL_u16_u16_600_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/MUL_u16_u16_600_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(335)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(335)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(335) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:MUL_u16_u16_600_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(335), ack => MUL_u16_u16_600_inst_req_1); -- 
    try1_cp_element_group_335: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_335"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(337) & try1_CP_1680_elements(340);
      gj_try1_cp_element_group_335 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(335), clk => clk, reset => reset); --
    end block;
    -- CP-element group 336:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	334 
    -- CP-element group 336: successors 
    -- CP-element group 336: marked-successors 
    -- CP-element group 336: 	323 
    -- CP-element group 336: 	327 
    -- CP-element group 336: 	334 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/MUL_u16_u16_600_sample_completed_
      -- CP-element group 336: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/MUL_u16_u16_600_Sample/$exit
      -- CP-element group 336: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/MUL_u16_u16_600_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(336)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(336)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(336) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:MUL_u16_u16_600_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_u16_u16_600_inst_ack_0, ack => try1_CP_1680_elements(336)); -- 
    -- CP-element group 337:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	335 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337: marked-successors 
    -- CP-element group 337: 	335 
    -- CP-element group 337:  members (3) 
      -- CP-element group 337: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/MUL_u16_u16_600_update_completed_
      -- CP-element group 337: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/MUL_u16_u16_600_Update/$exit
      -- CP-element group 337: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/MUL_u16_u16_600_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(337)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(337)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(337) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:MUL_u16_u16_600_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUL_u16_u16_600_inst_ack_1, ack => try1_CP_1680_elements(337)); -- 
    -- CP-element group 338:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	333 
    -- CP-element group 338: 	337 
    -- CP-element group 338: marked-predecessors 
    -- CP-element group 338: 	340 
    -- CP-element group 338: 	365 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	340 
    -- CP-element group 338:  members (9) 
      -- CP-element group 338: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_sample_start_
      -- CP-element group 338: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_Sample/$entry
      -- CP-element group 338: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_Sample/array_obj_ref_597_Split/$entry
      -- CP-element group 338: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_Sample/array_obj_ref_597_Split/$exit
      -- CP-element group 338: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_Sample/array_obj_ref_597_Split/split_req
      -- CP-element group 338: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_Sample/array_obj_ref_597_Split/split_ack
      -- CP-element group 338: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_Sample/word_access_start/$entry
      -- CP-element group 338: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_Sample/word_access_start/word_0/$entry
      -- CP-element group 338: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(338)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(338)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(338) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_597_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(338), ack => array_obj_ref_597_store_0_req_0); -- 
    try1_cp_element_group_338: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_338"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= try1_CP_1680_elements(333) & try1_CP_1680_elements(337) & try1_CP_1680_elements(340) & try1_CP_1680_elements(365);
      gj_try1_cp_element_group_338 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(338), clk => clk, reset => reset); --
    end block;
    -- CP-element group 339:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: marked-predecessors 
    -- CP-element group 339: 	341 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	341 
    -- CP-element group 339:  members (5) 
      -- CP-element group 339: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_update_start_
      -- CP-element group 339: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_Update/word_access_complete/$entry
      -- CP-element group 339: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_Update/word_access_complete/word_0/$entry
      -- CP-element group 339: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(339)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(339)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(339) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_597_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(339), ack => array_obj_ref_597_store_0_req_1); -- 
    try1_cp_element_group_339: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_339"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(341);
      gj_try1_cp_element_group_339 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(339), clk => clk, reset => reset); --
    end block;
    -- CP-element group 340:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	338 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	364 
    -- CP-element group 340: 	365 
    -- CP-element group 340: marked-successors 
    -- CP-element group 340: 	331 
    -- CP-element group 340: 	335 
    -- CP-element group 340: 	338 
    -- CP-element group 340:  members (5) 
      -- CP-element group 340: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_sample_completed_
      -- CP-element group 340: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_Sample/$exit
      -- CP-element group 340: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_Sample/word_access_start/$exit
      -- CP-element group 340: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_Sample/word_access_start/word_0/$exit
      -- CP-element group 340: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(340)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(340)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(340) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_597_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_597_store_0_ack_0, ack => try1_CP_1680_elements(340)); -- 
    -- CP-element group 341:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	339 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	366 
    -- CP-element group 341: marked-successors 
    -- CP-element group 341: 	339 
    -- CP-element group 341:  members (5) 
      -- CP-element group 341: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_update_completed_
      -- CP-element group 341: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_Update/$exit
      -- CP-element group 341: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_Update/word_access_complete/$exit
      -- CP-element group 341: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_Update/word_access_complete/word_0/$exit
      -- CP-element group 341: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(341)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(341)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(341) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_597_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_597_store_0_ack_1, ack => try1_CP_1680_elements(341)); -- 
    -- CP-element group 342:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	347 
    -- CP-element group 342: 	351 
    -- CP-element group 342: marked-predecessors 
    -- CP-element group 342: 	352 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	352 
    -- CP-element group 342:  members (3) 
      -- CP-element group 342: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u16_u16_606_sample_start_
      -- CP-element group 342: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u16_u16_606_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u16_u16_606_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(342)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(342)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(342) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u16_u16_606_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(342), ack => ADD_u16_u16_606_inst_req_0); -- 
    try1_cp_element_group_342: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_342"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(347) & try1_CP_1680_elements(351) & try1_CP_1680_elements(352);
      gj_try1_cp_element_group_342 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(342), clk => clk, reset => reset); --
    end block;
    -- CP-element group 343:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: marked-predecessors 
    -- CP-element group 343: 	353 
    -- CP-element group 343: 	356 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	353 
    -- CP-element group 343:  members (3) 
      -- CP-element group 343: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u16_u16_606_update_start_
      -- CP-element group 343: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u16_u16_606_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u16_u16_606_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(343)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(343)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(343) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u16_u16_606_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(343), ack => ADD_u16_u16_606_inst_req_1); -- 
    try1_cp_element_group_343: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_343"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(353) & try1_CP_1680_elements(356);
      gj_try1_cp_element_group_343 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(343), clk => clk, reset => reset); --
    end block;
    -- CP-element group 344:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	302 
    -- CP-element group 344: marked-predecessors 
    -- CP-element group 344: 	346 
    -- CP-element group 344: 	356 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	346 
    -- CP-element group 344:  members (5) 
      -- CP-element group 344: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_sample_start_
      -- CP-element group 344: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_Sample/$entry
      -- CP-element group 344: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_Sample/word_access_start/$entry
      -- CP-element group 344: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_Sample/word_access_start/word_0/$entry
      -- CP-element group 344: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(344)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(344)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(344) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_total_603_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(344), ack => LOAD_total_603_load_0_req_0); -- 
    try1_cp_element_group_344: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_344"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(302) & try1_CP_1680_elements(346) & try1_CP_1680_elements(356);
      gj_try1_cp_element_group_344 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(344), clk => clk, reset => reset); --
    end block;
    -- CP-element group 345:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: marked-predecessors 
    -- CP-element group 345: 	347 
    -- CP-element group 345: 	352 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	347 
    -- CP-element group 345:  members (5) 
      -- CP-element group 345: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_update_start_
      -- CP-element group 345: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_Update/word_access_complete/$entry
      -- CP-element group 345: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_Update/word_access_complete/word_0/$entry
      -- CP-element group 345: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(345)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(345)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(345) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_total_603_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(345), ack => LOAD_total_603_load_0_req_1); -- 
    try1_cp_element_group_345: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_345"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(347) & try1_CP_1680_elements(352);
      gj_try1_cp_element_group_345 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(345), clk => clk, reset => reset); --
    end block;
    -- CP-element group 346:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	344 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	363 
    -- CP-element group 346: marked-successors 
    -- CP-element group 346: 	344 
    -- CP-element group 346:  members (5) 
      -- CP-element group 346: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_sample_completed_
      -- CP-element group 346: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_Sample/$exit
      -- CP-element group 346: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_Sample/word_access_start/$exit
      -- CP-element group 346: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_Sample/word_access_start/word_0/$exit
      -- CP-element group 346: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(346)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(346)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(346) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_total_603_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_total_603_load_0_ack_0, ack => try1_CP_1680_elements(346)); -- 
    -- CP-element group 347:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	345 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	342 
    -- CP-element group 347: marked-successors 
    -- CP-element group 347: 	345 
    -- CP-element group 347:  members (9) 
      -- CP-element group 347: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_update_completed_
      -- CP-element group 347: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_Update/$exit
      -- CP-element group 347: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_Update/word_access_complete/$exit
      -- CP-element group 347: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_Update/word_access_complete/word_0/$exit
      -- CP-element group 347: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_Update/word_access_complete/word_0/ca
      -- CP-element group 347: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_Update/LOAD_total_603_Merge/$entry
      -- CP-element group 347: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_Update/LOAD_total_603_Merge/$exit
      -- CP-element group 347: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_Update/LOAD_total_603_Merge/merge_req
      -- CP-element group 347: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_Update/LOAD_total_603_Merge/merge_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(347)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(347)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(347) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_total_603_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_total_603_load_0_ack_1, ack => try1_CP_1680_elements(347)); -- 
    -- CP-element group 348:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	308 
    -- CP-element group 348: 	364 
    -- CP-element group 348: marked-predecessors 
    -- CP-element group 348: 	350 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	350 
    -- CP-element group 348:  members (5) 
      -- CP-element group 348: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_sample_start_
      -- CP-element group 348: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_Sample/$entry
      -- CP-element group 348: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_Sample/word_access_start/$entry
      -- CP-element group 348: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_Sample/word_access_start/word_0/$entry
      -- CP-element group 348: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(348)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(348)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(348) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_605_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(348), ack => array_obj_ref_605_load_0_req_0); -- 
    try1_cp_element_group_348: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_348"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(308) & try1_CP_1680_elements(364) & try1_CP_1680_elements(350);
      gj_try1_cp_element_group_348 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(348), clk => clk, reset => reset); --
    end block;
    -- CP-element group 349:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: marked-predecessors 
    -- CP-element group 349: 	351 
    -- CP-element group 349: 	352 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	351 
    -- CP-element group 349:  members (5) 
      -- CP-element group 349: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_update_start_
      -- CP-element group 349: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_Update/$entry
      -- CP-element group 349: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_Update/word_access_complete/$entry
      -- CP-element group 349: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_Update/word_access_complete/word_0/$entry
      -- CP-element group 349: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(349)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(349)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(349) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_605_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(349), ack => array_obj_ref_605_load_0_req_1); -- 
    try1_cp_element_group_349: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_349"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(351) & try1_CP_1680_elements(352);
      gj_try1_cp_element_group_349 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(349), clk => clk, reset => reset); --
    end block;
    -- CP-element group 350:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	348 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	365 
    -- CP-element group 350: marked-successors 
    -- CP-element group 350: 	306 
    -- CP-element group 350: 	348 
    -- CP-element group 350:  members (5) 
      -- CP-element group 350: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_sample_completed_
      -- CP-element group 350: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_Sample/$exit
      -- CP-element group 350: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_Sample/word_access_start/$exit
      -- CP-element group 350: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_Sample/word_access_start/word_0/$exit
      -- CP-element group 350: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(350)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(350)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(350) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_605_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_605_load_0_ack_0, ack => try1_CP_1680_elements(350)); -- 
    -- CP-element group 351:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	349 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	342 
    -- CP-element group 351: marked-successors 
    -- CP-element group 351: 	349 
    -- CP-element group 351:  members (9) 
      -- CP-element group 351: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_update_completed_
      -- CP-element group 351: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_Update/$exit
      -- CP-element group 351: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_Update/word_access_complete/$exit
      -- CP-element group 351: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_Update/word_access_complete/word_0/$exit
      -- CP-element group 351: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_Update/word_access_complete/word_0/ca
      -- CP-element group 351: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_Update/array_obj_ref_605_Merge/$entry
      -- CP-element group 351: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_Update/array_obj_ref_605_Merge/$exit
      -- CP-element group 351: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_Update/array_obj_ref_605_Merge/merge_req
      -- CP-element group 351: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_605_Update/array_obj_ref_605_Merge/merge_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(351)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(351)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(351) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_605_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_605_load_0_ack_1, ack => try1_CP_1680_elements(351)); -- 
    -- CP-element group 352:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	342 
    -- CP-element group 352: successors 
    -- CP-element group 352: marked-successors 
    -- CP-element group 352: 	342 
    -- CP-element group 352: 	345 
    -- CP-element group 352: 	349 
    -- CP-element group 352:  members (3) 
      -- CP-element group 352: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u16_u16_606_sample_completed_
      -- CP-element group 352: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u16_u16_606_Sample/$exit
      -- CP-element group 352: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u16_u16_606_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(352)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(352)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(352) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u16_u16_606_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_606_inst_ack_0, ack => try1_CP_1680_elements(352)); -- 
    -- CP-element group 353:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	343 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	354 
    -- CP-element group 353: marked-successors 
    -- CP-element group 353: 	343 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u16_u16_606_update_completed_
      -- CP-element group 353: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u16_u16_606_Update/$exit
      -- CP-element group 353: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u16_u16_606_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(353)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(353)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(353) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u16_u16_606_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u16_u16_606_inst_ack_1, ack => try1_CP_1680_elements(353)); -- 
    -- CP-element group 354:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	302 
    -- CP-element group 354: 	353 
    -- CP-element group 354: 	363 
    -- CP-element group 354: marked-predecessors 
    -- CP-element group 354: 	356 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	356 
    -- CP-element group 354:  members (9) 
      -- CP-element group 354: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_sample_start_
      -- CP-element group 354: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_Sample/$entry
      -- CP-element group 354: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_Sample/STORE_total_602_Split/$entry
      -- CP-element group 354: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_Sample/STORE_total_602_Split/$exit
      -- CP-element group 354: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_Sample/STORE_total_602_Split/split_req
      -- CP-element group 354: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_Sample/STORE_total_602_Split/split_ack
      -- CP-element group 354: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_Sample/word_access_start/$entry
      -- CP-element group 354: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_Sample/word_access_start/word_0/$entry
      -- CP-element group 354: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(354)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(354)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(354) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:STORE_total_602_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(354), ack => STORE_total_602_store_0_req_0); -- 
    try1_cp_element_group_354: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_354"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= try1_CP_1680_elements(302) & try1_CP_1680_elements(353) & try1_CP_1680_elements(363) & try1_CP_1680_elements(356);
      gj_try1_cp_element_group_354 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(354), clk => clk, reset => reset); --
    end block;
    -- CP-element group 355:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: marked-predecessors 
    -- CP-element group 355: 	357 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	357 
    -- CP-element group 355:  members (5) 
      -- CP-element group 355: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_update_start_
      -- CP-element group 355: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_Update/$entry
      -- CP-element group 355: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_Update/word_access_complete/$entry
      -- CP-element group 355: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_Update/word_access_complete/word_0/$entry
      -- CP-element group 355: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(355)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(355)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(355) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:STORE_total_602_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(355), ack => STORE_total_602_store_0_req_1); -- 
    try1_cp_element_group_355: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_355"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(357);
      gj_try1_cp_element_group_355 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(355), clk => clk, reset => reset); --
    end block;
    -- CP-element group 356:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	354 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	366 
    -- CP-element group 356: marked-successors 
    -- CP-element group 356: 	343 
    -- CP-element group 356: 	344 
    -- CP-element group 356: 	354 
    -- CP-element group 356:  members (6) 
      -- CP-element group 356: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_sample_completed_
      -- CP-element group 356: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_Sample/$exit
      -- CP-element group 356: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_Sample/word_access_start/$exit
      -- CP-element group 356: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_Sample/word_access_start/word_0/$exit
      -- CP-element group 356: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_Sample/word_access_start/word_0/ra
      -- CP-element group 356: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ring_reenable_memory_space_7
      -- 
    -- logger for CP element group try1_CP_1680_elements(356)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(356)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(356) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:STORE_total_602_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_total_602_store_0_ack_0, ack => try1_CP_1680_elements(356)); -- 
    -- CP-element group 357:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	355 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	366 
    -- CP-element group 357: marked-successors 
    -- CP-element group 357: 	355 
    -- CP-element group 357:  members (5) 
      -- CP-element group 357: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_update_completed_
      -- CP-element group 357: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_Update/$exit
      -- CP-element group 357: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_Update/word_access_complete/$exit
      -- CP-element group 357: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_Update/word_access_complete/word_0/$exit
      -- CP-element group 357: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/STORE_total_602_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(357)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(357)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(357) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:STORE_total_602_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_total_602_store_0_ack_1, ack => try1_CP_1680_elements(357)); -- 
    -- CP-element group 358:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	308 
    -- CP-element group 358: marked-predecessors 
    -- CP-element group 358: 	360 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	360 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u32_u32_611_sample_start_
      -- CP-element group 358: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u32_u32_611_Sample/$entry
      -- CP-element group 358: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u32_u32_611_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(358)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(358)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(358) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u32_u32_611_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(358), ack => ADD_u32_u32_611_inst_req_0); -- 
    try1_cp_element_group_358: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_358"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(308) & try1_CP_1680_elements(360);
      gj_try1_cp_element_group_358 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(358), clk => clk, reset => reset); --
    end block;
    -- CP-element group 359:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	307 
    -- CP-element group 359: marked-predecessors 
    -- CP-element group 359: 	361 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	361 
    -- CP-element group 359:  members (3) 
      -- CP-element group 359: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u32_u32_611_update_start_
      -- CP-element group 359: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u32_u32_611_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u32_u32_611_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(359)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(359)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(359) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u32_u32_611_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(359), ack => ADD_u32_u32_611_inst_req_1); -- 
    try1_cp_element_group_359: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_359"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(307) & try1_CP_1680_elements(361);
      gj_try1_cp_element_group_359 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(359), clk => clk, reset => reset); --
    end block;
    -- CP-element group 360:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	358 
    -- CP-element group 360: successors 
    -- CP-element group 360: marked-successors 
    -- CP-element group 360: 	306 
    -- CP-element group 360: 	358 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u32_u32_611_sample_completed_
      -- CP-element group 360: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u32_u32_611_Sample/$exit
      -- CP-element group 360: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u32_u32_611_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(360)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(360)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(360) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u32_u32_611_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_611_inst_ack_0, ack => try1_CP_1680_elements(360)); -- 
    -- CP-element group 361:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	359 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	303 
    -- CP-element group 361: marked-successors 
    -- CP-element group 361: 	305 
    -- CP-element group 361: 	359 
    -- CP-element group 361:  members (3) 
      -- CP-element group 361: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u32_u32_611_update_completed_
      -- CP-element group 361: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u32_u32_611_Update/$exit
      -- CP-element group 361: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ADD_u32_u32_611_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(361)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(361)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(361) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u32_u32_611_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_611_inst_ack_1, ack => try1_CP_1680_elements(361)); -- 
    -- CP-element group 362:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	302 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	303 
    -- CP-element group 362:  members (1) 
      -- CP-element group 362: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group try1_CP_1680_elements(362)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(362)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(362) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(362) is a control-delay.
    cp_element_362_delay: control_delay_element  generic map(name => " 362_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(302), ack => try1_CP_1680_elements(362), clk => clk, reset =>reset);
    -- CP-element group 363:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	346 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	354 
    -- CP-element group 363:  members (1) 
      -- CP-element group 363: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/LOAD_total_603_STORE_total_602_delay
      -- 
    -- logger for CP element group try1_CP_1680_elements(363)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(363)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(363) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(363) is a control-delay.
    cp_element_363_delay: control_delay_element  generic map(name => " 363_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(346), ack => try1_CP_1680_elements(363), clk => clk, reset =>reset);
    -- CP-element group 364:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	340 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	348 
    -- CP-element group 364:  members (1) 
      -- CP-element group 364: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/array_obj_ref_597_array_obj_ref_605_delay
      -- 
    -- logger for CP element group try1_CP_1680_elements(364)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(364)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(364) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(364) is a control-delay.
    cp_element_364_delay: control_delay_element  generic map(name => " 364_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(340), ack => try1_CP_1680_elements(364), clk => clk, reset =>reset);
    -- CP-element group 365:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	340 
    -- CP-element group 365: 	350 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365: marked-successors 
    -- CP-element group 365: 	338 
    -- CP-element group 365:  members (1) 
      -- CP-element group 365: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/ring_reenable_memory_space_2
      -- 
    -- logger for CP element group try1_CP_1680_elements(365)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(365)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(365) fired."); 
        -- 
      end if; --
    end process; 
    try1_cp_element_group_365: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_365"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(340) & try1_CP_1680_elements(350);
      gj_try1_cp_element_group_365 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(365), clk => clk, reset => reset); --
    end block;
    -- CP-element group 366:  join  transition  bypass  pipeline-parent 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	341 
    -- CP-element group 366: 	356 
    -- CP-element group 366: 	357 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	299 
    -- CP-element group 366:  members (1) 
      -- CP-element group 366: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/do_while_stmt_577_loop_body/$exit
      -- 
    -- logger for CP element group try1_CP_1680_elements(366)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(366)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(366) fired."); 
        -- 
      end if; --
    end process; 
    try1_cp_element_group_366: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 7,2 => 7,3 => 7);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_366"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= try1_CP_1680_elements(341) & try1_CP_1680_elements(356) & try1_CP_1680_elements(357) & try1_CP_1680_elements(365);
      gj_try1_cp_element_group_366 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(366), clk => clk, reset => reset); --
    end block;
    -- CP-element group 367:  transition  input  bypass  pipeline-parent 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	298 
    -- CP-element group 367: successors 
    -- CP-element group 367:  members (2) 
      -- CP-element group 367: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/loop_exit/$exit
      -- CP-element group 367: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/loop_exit/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(367)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(367)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(367) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:do_while_stmt_577_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_577_branch_ack_0, ack => try1_CP_1680_elements(367)); -- 
    -- CP-element group 368:  transition  input  bypass  pipeline-parent 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	298 
    -- CP-element group 368: successors 
    -- CP-element group 368:  members (2) 
      -- CP-element group 368: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/loop_taken/$exit
      -- CP-element group 368: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/loop_taken/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(368)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(368)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(368) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:do_while_stmt_577_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_577_branch_ack_1, ack => try1_CP_1680_elements(368)); -- 
    -- CP-element group 369:  transition  bypass  pipeline-parent 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	296 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	294 
    -- CP-element group 369:  members (1) 
      -- CP-element group 369: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_576/do_while_stmt_577/$exit
      -- 
    -- logger for CP element group try1_CP_1680_elements(369)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(369)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(369) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(369) <= try1_CP_1680_elements(296);
    -- CP-element group 370:  join  transition  output  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	372 
    -- CP-element group 370: 	374 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	375 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/call_stmt_624_sample_start_
      -- CP-element group 370: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/call_stmt_624_Sample/$entry
      -- CP-element group 370: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/call_stmt_624_Sample/crr
      -- 
    -- logger for CP element group try1_CP_1680_elements(370)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(370)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(370) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:call_stmt_624_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_3779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(370), ack => call_stmt_624_call_req_0); -- 
    try1_cp_element_group_370: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_370"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(372) & try1_CP_1680_elements(374);
      gj_try1_cp_element_group_370 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(370), clk => clk, reset => reset); --
    end block;
    -- CP-element group 371:  transition  input  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	294 
    -- CP-element group 371: successors 
    -- CP-element group 371:  members (3) 
      -- CP-element group 371: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/ADD_u12_u12_621_sample_completed_
      -- CP-element group 371: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/ADD_u12_u12_621_Sample/$exit
      -- CP-element group 371: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/ADD_u12_u12_621_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(371)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(371)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(371) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_621_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_621_inst_ack_0, ack => try1_CP_1680_elements(371)); -- 
    -- CP-element group 372:  transition  input  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	294 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	370 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/ADD_u12_u12_621_update_completed_
      -- CP-element group 372: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/ADD_u12_u12_621_Update/$exit
      -- CP-element group 372: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/ADD_u12_u12_621_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(372)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(372)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(372) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_621_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_621_inst_ack_1, ack => try1_CP_1680_elements(372)); -- 
    -- CP-element group 373:  transition  input  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	294 
    -- CP-element group 373: successors 
    -- CP-element group 373:  members (5) 
      -- CP-element group 373: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_sample_completed_
      -- CP-element group 373: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_Sample/$exit
      -- CP-element group 373: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_Sample/word_access_start/$exit
      -- CP-element group 373: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_Sample/word_access_start/word_0/$exit
      -- CP-element group 373: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(373)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(373)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(373) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_total_622_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_total_622_load_0_ack_0, ack => try1_CP_1680_elements(373)); -- 
    -- CP-element group 374:  transition  input  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	294 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	370 
    -- CP-element group 374:  members (9) 
      -- CP-element group 374: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_update_completed_
      -- CP-element group 374: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_Update/$exit
      -- CP-element group 374: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_Update/word_access_complete/$exit
      -- CP-element group 374: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_Update/word_access_complete/word_0/$exit
      -- CP-element group 374: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_Update/word_access_complete/word_0/ca
      -- CP-element group 374: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_Update/LOAD_total_622_Merge/$entry
      -- CP-element group 374: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_Update/LOAD_total_622_Merge/$exit
      -- CP-element group 374: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_Update/LOAD_total_622_Merge/merge_req
      -- CP-element group 374: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_total_622_Update/LOAD_total_622_Merge/merge_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(374)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(374)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(374) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_total_622_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_total_622_load_0_ack_1, ack => try1_CP_1680_elements(374)); -- 
    -- CP-element group 375:  transition  input  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	370 
    -- CP-element group 375: successors 
    -- CP-element group 375:  members (3) 
      -- CP-element group 375: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/call_stmt_624_sample_completed_
      -- CP-element group 375: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/call_stmt_624_Sample/$exit
      -- CP-element group 375: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/call_stmt_624_Sample/cra
      -- 
    -- logger for CP element group try1_CP_1680_elements(375)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(375)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(375) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:call_stmt_624_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_3780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_624_call_ack_0, ack => try1_CP_1680_elements(375)); -- 
    -- CP-element group 376:  transition  input  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	294 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	388 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/call_stmt_624_update_completed_
      -- CP-element group 376: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/call_stmt_624_Update/$exit
      -- CP-element group 376: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/call_stmt_624_Update/cca
      -- 
    -- logger for CP element group try1_CP_1680_elements(376)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(376)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(376) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:call_stmt_624_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_3785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_624_call_ack_1, ack => try1_CP_1680_elements(376)); -- 
    -- CP-element group 377:  transition  input  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	294 
    -- CP-element group 377: successors 
    -- CP-element group 377:  members (5) 
      -- CP-element group 377: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_sample_completed_
      -- CP-element group 377: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_Sample/$exit
      -- CP-element group 377: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_Sample/word_access_start/$exit
      -- CP-element group 377: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_Sample/word_access_start/word_0/$exit
      -- CP-element group 377: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(377)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(377)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(377) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_zer_626_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_zer_626_load_0_ack_0, ack => try1_CP_1680_elements(377)); -- 
    -- CP-element group 378:  transition  input  output  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	294 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	379 
    -- CP-element group 378:  members (12) 
      -- CP-element group 378: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/CONCAT_u4_u16_630_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_update_completed_
      -- CP-element group 378: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_Update/$exit
      -- CP-element group 378: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_Update/word_access_complete/$exit
      -- CP-element group 378: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_Update/word_access_complete/word_0/$exit
      -- CP-element group 378: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_Update/word_access_complete/word_0/ca
      -- CP-element group 378: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_Update/LOAD_zer_626_Merge/$entry
      -- CP-element group 378: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_Update/LOAD_zer_626_Merge/$exit
      -- CP-element group 378: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_Update/LOAD_zer_626_Merge/merge_req
      -- CP-element group 378: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/LOAD_zer_626_Update/LOAD_zer_626_Merge/merge_ack
      -- CP-element group 378: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/CONCAT_u4_u16_630_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/CONCAT_u4_u16_630_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(378)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(378)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(378) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:LOAD_zer_626_load_0_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:CONCAT_u4_u16_630_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_3817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_zer_626_load_0_ack_1, ack => try1_CP_1680_elements(378)); -- 
    rr_3826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(378), ack => CONCAT_u4_u16_630_inst_req_0); -- 
    -- CP-element group 379:  transition  input  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	378 
    -- CP-element group 379: successors 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/CONCAT_u4_u16_630_sample_completed_
      -- CP-element group 379: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/CONCAT_u4_u16_630_Sample/$exit
      -- CP-element group 379: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/CONCAT_u4_u16_630_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(379)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(379)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(379) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:CONCAT_u4_u16_630_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u4_u16_630_inst_ack_0, ack => try1_CP_1680_elements(379)); -- 
    -- CP-element group 380:  fork  transition  input  output  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	294 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	383 
    -- CP-element group 380: 	381 
    -- CP-element group 380:  members (32) 
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/CONCAT_u4_u16_630_update_completed_
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/CONCAT_u4_u16_630_Update/$exit
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/CONCAT_u4_u16_630_Update/ca
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_add_632_sample_start_
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_add_632_Sample/$entry
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_add_632_Sample/req
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_word_address_calculated
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_root_address_calculated
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_offset_calculated
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_index_resized_0
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_index_scaled_0
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_index_computed_0
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_index_resize_0/$entry
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_index_resize_0/$exit
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_index_resize_0/index_resize_req
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_index_resize_0/index_resize_ack
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_index_scale_0/$entry
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_index_scale_0/$exit
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_index_scale_0/scale_rename_req
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_index_scale_0/scale_rename_ack
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_final_index_sum_regn/$entry
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_final_index_sum_regn/$exit
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_final_index_sum_regn/req
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_final_index_sum_regn/ack
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_base_plus_offset/$entry
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_base_plus_offset/$exit
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_base_plus_offset/sum_rename_req
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_base_plus_offset/sum_rename_ack
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_word_addrgen/$entry
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_word_addrgen/$exit
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_word_addrgen/root_register_req
      -- CP-element group 380: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(380)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(380)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(380) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:CONCAT_u4_u16_630_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:WPIPE_acc_mem_add_632_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_3832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u4_u16_630_inst_ack_1, ack => try1_CP_1680_elements(380)); -- 
    req_3840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(380), ack => WPIPE_acc_mem_add_632_inst_req_0); -- 
    -- CP-element group 381:  transition  input  output  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	380 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	382 
    -- CP-element group 381:  members (6) 
      -- CP-element group 381: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_add_632_sample_completed_
      -- CP-element group 381: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_add_632_update_start_
      -- CP-element group 381: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_add_632_Sample/$exit
      -- CP-element group 381: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_add_632_Sample/ack
      -- CP-element group 381: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_add_632_Update/$entry
      -- CP-element group 381: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_add_632_Update/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(381)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(381)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(381) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:WPIPE_acc_mem_add_632_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:WPIPE_acc_mem_add_632_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_acc_mem_add_632_inst_ack_0, ack => try1_CP_1680_elements(381)); -- 
    req_3845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(381), ack => WPIPE_acc_mem_add_632_inst_req_1); -- 
    -- CP-element group 382:  transition  input  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	381 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	389 
    -- CP-element group 382:  members (3) 
      -- CP-element group 382: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_add_632_update_completed_
      -- CP-element group 382: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_add_632_Update/$exit
      -- CP-element group 382: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_add_632_Update/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(382)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(382)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(382) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:WPIPE_acc_mem_add_632_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_acc_mem_add_632_inst_ack_1, ack => try1_CP_1680_elements(382)); -- 
    -- CP-element group 383:  join  transition  output  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	388 
    -- CP-element group 383: 	380 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	384 
    -- CP-element group 383:  members (5) 
      -- CP-element group 383: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_sample_start_
      -- CP-element group 383: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_Sample/$entry
      -- CP-element group 383: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_Sample/word_access_start/$entry
      -- CP-element group 383: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_Sample/word_access_start/word_0/$entry
      -- CP-element group 383: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(383)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(383)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(383) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_637_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(383), ack => array_obj_ref_637_load_0_req_0); -- 
    try1_cp_element_group_383: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_383"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(388) & try1_CP_1680_elements(380);
      gj_try1_cp_element_group_383 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(383), clk => clk, reset => reset); --
    end block;
    -- CP-element group 384:  transition  input  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	383 
    -- CP-element group 384: successors 
    -- CP-element group 384:  members (5) 
      -- CP-element group 384: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_sample_completed_
      -- CP-element group 384: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_Sample/$exit
      -- CP-element group 384: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_Sample/word_access_start/$exit
      -- CP-element group 384: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_Sample/word_access_start/word_0/$exit
      -- CP-element group 384: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(384)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(384)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(384) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_637_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_637_load_0_ack_0, ack => try1_CP_1680_elements(384)); -- 
    -- CP-element group 385:  transition  input  output  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	294 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	386 
    -- CP-element group 385:  members (12) 
      -- CP-element group 385: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_update_completed_
      -- CP-element group 385: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_Update/$exit
      -- CP-element group 385: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_Update/word_access_complete/$exit
      -- CP-element group 385: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_Update/word_access_complete/word_0/$exit
      -- CP-element group 385: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_Update/word_access_complete/word_0/ca
      -- CP-element group 385: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_Update/array_obj_ref_637_Merge/$entry
      -- CP-element group 385: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_Update/array_obj_ref_637_Merge/$exit
      -- CP-element group 385: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_Update/array_obj_ref_637_Merge/merge_req
      -- CP-element group 385: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/array_obj_ref_637_Update/array_obj_ref_637_Merge/merge_ack
      -- CP-element group 385: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_635_sample_start_
      -- CP-element group 385: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_635_Sample/$entry
      -- CP-element group 385: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_635_Sample/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(385)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(385)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(385) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_637_load_0_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:WPIPE_acc_mem_635_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_3904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_637_load_0_ack_1, ack => try1_CP_1680_elements(385)); -- 
    req_3917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(385), ack => WPIPE_acc_mem_635_inst_req_0); -- 
    -- CP-element group 386:  transition  input  output  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	385 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	387 
    -- CP-element group 386:  members (6) 
      -- CP-element group 386: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_635_sample_completed_
      -- CP-element group 386: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_635_update_start_
      -- CP-element group 386: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_635_Sample/$exit
      -- CP-element group 386: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_635_Sample/ack
      -- CP-element group 386: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_635_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_635_Update/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(386)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(386)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(386) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:WPIPE_acc_mem_635_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:WPIPE_acc_mem_635_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_acc_mem_635_inst_ack_0, ack => try1_CP_1680_elements(386)); -- 
    req_3922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(386), ack => WPIPE_acc_mem_635_inst_req_1); -- 
    -- CP-element group 387:  transition  input  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	386 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	389 
    -- CP-element group 387:  members (3) 
      -- CP-element group 387: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_635_update_completed_
      -- CP-element group 387: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_635_Update/$exit
      -- CP-element group 387: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/WPIPE_acc_mem_635_Update/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(387)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(387)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(387) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:WPIPE_acc_mem_635_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_acc_mem_635_inst_ack_1, ack => try1_CP_1680_elements(387)); -- 
    -- CP-element group 388:  transition  delay-element  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	376 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	383 
    -- CP-element group 388:  members (1) 
      -- CP-element group 388: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/call_stmt_624_array_obj_ref_637_delay
      -- 
    -- logger for CP element group try1_CP_1680_elements(388)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(388)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(388) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(388) is a control-delay.
    cp_element_388_delay: control_delay_element  generic map(name => " 388_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(376), ack => try1_CP_1680_elements(388), clk => clk, reset =>reset);
    -- CP-element group 389:  join  transition  place  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	387 
    -- CP-element group 389: 	382 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	391 
    -- CP-element group 389:  members (6) 
      -- CP-element group 389: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638__exit__
      -- CP-element group 389: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639__entry__
      -- CP-element group 389: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/$entry
      -- CP-element group 389: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640__entry__
      -- CP-element group 389: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/branch_block_stmt_639__entry__
      -- CP-element group 389: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_624_to_assign_stmt_638/$exit
      -- 
    -- logger for CP element group try1_CP_1680_elements(389)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(389)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(389) fired."); 
        -- 
      end if; --
    end process; 
    try1_cp_element_group_389: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_389"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(387) & try1_CP_1680_elements(382);
      gj_try1_cp_element_group_389 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(389), clk => clk, reset => reset); --
    end block;
    -- CP-element group 390:  fork  transition  place  output  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	479 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	480 
    -- CP-element group 390: 	481 
    -- CP-element group 390: 	483 
    -- CP-element group 390: 	485 
    -- CP-element group 390: 	486 
    -- CP-element group 390: 	493 
    -- CP-element group 390: 	495 
    -- CP-element group 390: 	496 
    -- CP-element group 390: 	498 
    -- CP-element group 390: 	500 
    -- CP-element group 390: 	501 
    -- CP-element group 390: 	503 
    -- CP-element group 390: 	504 
    -- CP-element group 390: 	505 
    -- CP-element group 390: 	490 
    -- CP-element group 390: 	491 
    -- CP-element group 390: 	488 
    -- CP-element group 390:  members (61) 
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639__exit__
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730__entry__
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/$exit
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640__exit__
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/branch_block_stmt_639__exit__
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/$entry
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/call_stmt_705_update_start_
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_702_sample_start_
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_702_update_start_
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_702_Sample/$entry
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_702_Sample/rr
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_702_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_702_Update/cr
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/call_stmt_705_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/call_stmt_705_Update/ccr
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_709_update_start_
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_709_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_709_Update/cr
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_update_start_
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_word_address_calculated
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_root_address_calculated
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_Update/word_access_complete/$entry
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_Update/word_access_complete/word_0/$entry
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_Update/word_access_complete/word_0/cr
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_714_update_start_
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_714_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_714_Update/cr
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_update_start_
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_word_address_calculated
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_root_address_calculated
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_Update/word_access_complete/$entry
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_Update/word_access_complete/word_0/$entry
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_Update/word_access_complete/word_0/cr
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_719_update_start_
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_719_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_719_Update/cr
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_update_start_
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_word_address_calculated
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_root_address_calculated
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_Update/word_access_complete/$entry
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_Update/word_access_complete/word_0/$entry
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_Update/word_access_complete/word_0/cr
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_724_update_start_
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_724_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_724_Update/cr
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_update_start_
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_word_address_calculated
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_root_address_calculated
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_Update/word_access_complete/$entry
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_Update/word_access_complete/word_0/$entry
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_Update/word_access_complete/word_0/cr
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_729_sample_start_
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_729_update_start_
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_729_Sample/$entry
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_729_Sample/rr
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_729_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_729_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(390)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(390)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(390) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_702_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_702_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:call_stmt_705_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_709_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_707_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_714_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_712_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_719_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_717_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_724_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_722_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_729_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_729_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    rr_4499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(390), ack => ADD_u12_u12_702_inst_req_0); -- 
    cr_4504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(390), ack => ADD_u12_u12_702_inst_req_1); -- 
    ccr_4514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(390), ack => call_stmt_705_call_req_1); -- 
    cr_4528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(390), ack => slice_709_inst_req_1); -- 
    cr_4561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(390), ack => array_obj_ref_707_store_0_req_1); -- 
    cr_4575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(390), ack => slice_714_inst_req_1); -- 
    cr_4608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(390), ack => array_obj_ref_712_store_0_req_1); -- 
    cr_4622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(390), ack => slice_719_inst_req_1); -- 
    cr_4655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(390), ack => array_obj_ref_717_store_0_req_1); -- 
    cr_4669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(390), ack => slice_724_inst_req_1); -- 
    cr_4702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(390), ack => array_obj_ref_722_store_0_req_1); -- 
    rr_4711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(390), ack => ADD_u12_u12_729_inst_req_0); -- 
    cr_4716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(390), ack => ADD_u12_u12_729_inst_req_1); -- 
    try1_CP_1680_elements(390) <= try1_CP_1680_elements(479);
    -- CP-element group 391:  transition  place  bypass  pipeline-parent 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	389 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	397 
    -- CP-element group 391:  members (2) 
      -- CP-element group 391: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/$entry
      -- CP-element group 391: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640__entry__
      -- 
    -- logger for CP element group try1_CP_1680_elements(391)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(391)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(391) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(391) <= try1_CP_1680_elements(389);
    -- CP-element group 392:  merge  place  bypass  pipeline-parent 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	479 
    -- CP-element group 392:  members (1) 
      -- CP-element group 392: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640__exit__
      -- 
    -- logger for CP element group try1_CP_1680_elements(392)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(392)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(392) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(392) is bound as output of CP function.
    -- CP-element group 393:  merge  place  bypass  pipeline-parent 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	396 
    -- CP-element group 393:  members (1) 
      -- CP-element group 393: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/loop_back
      -- 
    -- logger for CP element group try1_CP_1680_elements(393)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(393)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(393) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(393) is bound as output of CP function.
    -- CP-element group 394:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	399 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	477 
    -- CP-element group 394: 	478 
    -- CP-element group 394:  members (3) 
      -- CP-element group 394: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/condition_done
      -- CP-element group 394: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/loop_exit/$entry
      -- CP-element group 394: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/loop_taken/$entry
      -- 
    -- logger for CP element group try1_CP_1680_elements(394)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(394)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(394) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(394) <= try1_CP_1680_elements(399);
    -- CP-element group 395:  branch  place  bypass  pipeline-parent 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	476 
    -- CP-element group 395: successors 
    -- CP-element group 395:  members (1) 
      -- CP-element group 395: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/loop_body_done
      -- 
    -- logger for CP element group try1_CP_1680_elements(395)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(395)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(395) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(395) <= try1_CP_1680_elements(476);
    -- CP-element group 396:  transition  bypass  pipeline-parent 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	393 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	405 
    -- CP-element group 396:  members (1) 
      -- CP-element group 396: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group try1_CP_1680_elements(396)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(396)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(396) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(396) <= try1_CP_1680_elements(393);
    -- CP-element group 397:  transition  bypass  pipeline-parent 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	391 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	407 
    -- CP-element group 397:  members (1) 
      -- CP-element group 397: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group try1_CP_1680_elements(397)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(397)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(397) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(397) <= try1_CP_1680_elements(391);
    -- CP-element group 398:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	470 
    -- CP-element group 398: 	401 
    -- CP-element group 398: 	402 
    -- CP-element group 398:  members (2) 
      -- CP-element group 398: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/$entry
      -- CP-element group 398: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/loop_body_start
      -- 
    -- logger for CP element group try1_CP_1680_elements(398)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(398)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(398) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(398) is bound as output of CP function.
    -- CP-element group 399:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	469 
    -- CP-element group 399: 	470 
    -- CP-element group 399: 	404 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	394 
    -- CP-element group 399:  members (1) 
      -- CP-element group 399: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/condition_evaluated
      -- 
    -- logger for CP element group try1_CP_1680_elements(399)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(399)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(399) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:do_while_stmt_640_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_3946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(399), ack => do_while_stmt_640_branch_req_0); -- 
    try1_cp_element_group_399: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_399"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(469) & try1_CP_1680_elements(470) & try1_CP_1680_elements(404);
      gj_try1_cp_element_group_399 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(399), clk => clk, reset => reset); --
    end block;
    -- CP-element group 400:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	401 
    -- CP-element group 400: marked-predecessors 
    -- CP-element group 400: 	404 
    -- CP-element group 400: successors 
    -- CP-element group 400:  members (2) 
      -- CP-element group 400: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/phi_stmt_642_sample_start__ps
      -- CP-element group 400: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/aggregated_phi_sample_req
      -- 
    -- logger for CP element group try1_CP_1680_elements(400)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(400)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(400) fired."); 
        -- 
      end if; --
    end process; 
    try1_cp_element_group_400: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_400"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(401) & try1_CP_1680_elements(404);
      gj_try1_cp_element_group_400 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(400), clk => clk, reset => reset); --
    end block;
    -- CP-element group 401:  join  transition  bypass  pipeline-parent 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	398 
    -- CP-element group 401: marked-predecessors 
    -- CP-element group 401: 	469 
    -- CP-element group 401: 	403 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	400 
    -- CP-element group 401:  members (1) 
      -- CP-element group 401: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/phi_stmt_642_sample_start_
      -- 
    -- logger for CP element group try1_CP_1680_elements(401)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(401)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(401) fired."); 
        -- 
      end if; --
    end process; 
    try1_cp_element_group_401: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_401"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(398) & try1_CP_1680_elements(469) & try1_CP_1680_elements(403);
      gj_try1_cp_element_group_401 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(401), clk => clk, reset => reset); --
    end block;
    -- CP-element group 402:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	398 
    -- CP-element group 402: marked-predecessors 
    -- CP-element group 402: 	468 
    -- CP-element group 402: 	452 
    -- CP-element group 402: 	404 
    -- CP-element group 402: 	420 
    -- CP-element group 402: 	424 
    -- CP-element group 402: 	436 
    -- CP-element group 402: successors 
    -- CP-element group 402:  members (3) 
      -- CP-element group 402: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/aggregated_phi_update_req
      -- CP-element group 402: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/phi_stmt_642_update_start__ps
      -- CP-element group 402: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/phi_stmt_642_update_start_
      -- 
    -- logger for CP element group try1_CP_1680_elements(402)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(402)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(402) fired."); 
        -- 
      end if; --
    end process; 
    try1_cp_element_group_402: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_402"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= try1_CP_1680_elements(398) & try1_CP_1680_elements(468) & try1_CP_1680_elements(452) & try1_CP_1680_elements(404) & try1_CP_1680_elements(420) & try1_CP_1680_elements(424) & try1_CP_1680_elements(436);
      gj_try1_cp_element_group_402 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(402), clk => clk, reset => reset); --
    end block;
    -- CP-element group 403:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	467 
    -- CP-element group 403: marked-successors 
    -- CP-element group 403: 	401 
    -- CP-element group 403:  members (3) 
      -- CP-element group 403: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/aggregated_phi_sample_ack
      -- CP-element group 403: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/phi_stmt_642_sample_completed_
      -- CP-element group 403: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/phi_stmt_642_sample_completed__ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(403)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(403)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(403) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(403) is bound as output of CP function.
    -- CP-element group 404:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	450 
    -- CP-element group 404: 	418 
    -- CP-element group 404: 	422 
    -- CP-element group 404: 	466 
    -- CP-element group 404: 	399 
    -- CP-element group 404: 	434 
    -- CP-element group 404: marked-successors 
    -- CP-element group 404: 	400 
    -- CP-element group 404: 	402 
    -- CP-element group 404:  members (3) 
      -- CP-element group 404: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/phi_stmt_642_update_completed__ps
      -- CP-element group 404: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/aggregated_phi_update_ack
      -- CP-element group 404: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/phi_stmt_642_update_completed_
      -- 
    -- logger for CP element group try1_CP_1680_elements(404)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(404)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(404) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(404) is bound as output of CP function.
    -- CP-element group 405:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	396 
    -- CP-element group 405: successors 
    -- CP-element group 405:  members (1) 
      -- CP-element group 405: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/phi_stmt_642_loopback_trigger
      -- 
    -- logger for CP element group try1_CP_1680_elements(405)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(405)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(405) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(405) <= try1_CP_1680_elements(396);
    -- CP-element group 406:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: successors 
    -- CP-element group 406:  members (2) 
      -- CP-element group 406: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/phi_stmt_642_loopback_sample_req_ps
      -- CP-element group 406: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/phi_stmt_642_loopback_sample_req
      -- 
    -- logger for CP element group try1_CP_1680_elements(406)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(406)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(406) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:phi_stmt_642_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_642_loopback_sample_req_3961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_642_loopback_sample_req_3961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(406), ack => phi_stmt_642_req_1); -- 
    -- Element group try1_CP_1680_elements(406) is bound as output of CP function.
    -- CP-element group 407:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	397 
    -- CP-element group 407: successors 
    -- CP-element group 407:  members (1) 
      -- CP-element group 407: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/phi_stmt_642_entry_trigger
      -- 
    -- logger for CP element group try1_CP_1680_elements(407)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(407)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(407) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(407) <= try1_CP_1680_elements(397);
    -- CP-element group 408:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: successors 
    -- CP-element group 408:  members (2) 
      -- CP-element group 408: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/phi_stmt_642_entry_sample_req_ps
      -- CP-element group 408: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/phi_stmt_642_entry_sample_req
      -- 
    -- logger for CP element group try1_CP_1680_elements(408)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(408)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(408) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:phi_stmt_642_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_642_entry_sample_req_3964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_642_entry_sample_req_3964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(408), ack => phi_stmt_642_req_0); -- 
    -- Element group try1_CP_1680_elements(408) is bound as output of CP function.
    -- CP-element group 409:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: successors 
    -- CP-element group 409:  members (2) 
      -- CP-element group 409: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/phi_stmt_642_phi_mux_ack
      -- CP-element group 409: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/phi_stmt_642_phi_mux_ack_ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(409)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(409)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(409) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:phi_stmt_642_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_642_phi_mux_ack_3967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 409_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_642_ack_0, ack => try1_CP_1680_elements(409)); -- 
    -- CP-element group 410:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: successors 
    -- CP-element group 410:  members (4) 
      -- CP-element group 410: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/type_cast_645_sample_start__ps
      -- CP-element group 410: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/type_cast_645_sample_completed__ps
      -- CP-element group 410: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/type_cast_645_sample_completed_
      -- CP-element group 410: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/type_cast_645_sample_start_
      -- 
    -- logger for CP element group try1_CP_1680_elements(410)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(410)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(410) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(410) is bound as output of CP function.
    -- CP-element group 411:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	413 
    -- CP-element group 411:  members (2) 
      -- CP-element group 411: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/type_cast_645_update_start_
      -- CP-element group 411: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/type_cast_645_update_start__ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(411)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(411)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(411) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(411) is bound as output of CP function.
    -- CP-element group 412:  join  transition  bypass  pipeline-parent 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	413 
    -- CP-element group 412: successors 
    -- CP-element group 412:  members (1) 
      -- CP-element group 412: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/type_cast_645_update_completed__ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(412)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(412)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(412) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(412) <= try1_CP_1680_elements(413);
    -- CP-element group 413:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	411 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	412 
    -- CP-element group 413:  members (1) 
      -- CP-element group 413: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/type_cast_645_update_completed_
      -- 
    -- logger for CP element group try1_CP_1680_elements(413)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(413)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(413) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(413) is a control-delay.
    cp_element_413_delay: control_delay_element  generic map(name => " 413_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(411), ack => try1_CP_1680_elements(413), clk => clk, reset =>reset);
    -- CP-element group 414:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	416 
    -- CP-element group 414:  members (4) 
      -- CP-element group 414: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/R_NH_646_Sample/req
      -- CP-element group 414: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/R_NH_646_Sample/$entry
      -- CP-element group 414: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/R_NH_646_sample_start_
      -- CP-element group 414: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/R_NH_646_sample_start__ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(414)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(414)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(414) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NH_691_646_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(414), ack => NH_691_646_buf_req_0); -- 
    -- Element group try1_CP_1680_elements(414) is bound as output of CP function.
    -- CP-element group 415:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	417 
    -- CP-element group 415:  members (4) 
      -- CP-element group 415: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/R_NH_646_Update/req
      -- CP-element group 415: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/R_NH_646_Update/$entry
      -- CP-element group 415: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/R_NH_646_update_start_
      -- CP-element group 415: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/R_NH_646_update_start__ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(415)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(415)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(415) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NH_691_646_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(415), ack => NH_691_646_buf_req_1); -- 
    -- Element group try1_CP_1680_elements(415) is bound as output of CP function.
    -- CP-element group 416:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	414 
    -- CP-element group 416: successors 
    -- CP-element group 416:  members (4) 
      -- CP-element group 416: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/R_NH_646_Sample/ack
      -- CP-element group 416: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/R_NH_646_Sample/$exit
      -- CP-element group 416: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/R_NH_646_sample_completed_
      -- CP-element group 416: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/R_NH_646_sample_completed__ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(416)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(416)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(416) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NH_691_646_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NH_691_646_buf_ack_0, ack => try1_CP_1680_elements(416)); -- 
    -- CP-element group 417:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	415 
    -- CP-element group 417: successors 
    -- CP-element group 417:  members (4) 
      -- CP-element group 417: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/R_NH_646_Update/ack
      -- CP-element group 417: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/R_NH_646_Update/$exit
      -- CP-element group 417: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/R_NH_646_update_completed_
      -- CP-element group 417: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/R_NH_646_update_completed__ps
      -- 
    -- logger for CP element group try1_CP_1680_elements(417)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(417)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(417) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NH_691_646_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NH_691_646_buf_ack_1, ack => try1_CP_1680_elements(417)); -- 
    -- CP-element group 418:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	404 
    -- CP-element group 418: marked-predecessors 
    -- CP-element group 418: 	420 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	420 
    -- CP-element group 418:  members (3) 
      -- CP-element group 418: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_651_Sample/rr
      -- CP-element group 418: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_651_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_651_sample_start_
      -- 
    -- logger for CP element group try1_CP_1680_elements(418)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(418)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(418) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_651_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(418), ack => ADD_u12_u12_651_inst_req_0); -- 
    try1_cp_element_group_418: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_418"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(404) & try1_CP_1680_elements(420);
      gj_try1_cp_element_group_418 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(418), clk => clk, reset => reset); --
    end block;
    -- CP-element group 419:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: marked-predecessors 
    -- CP-element group 419: 	421 
    -- CP-element group 419: 	440 
    -- CP-element group 419: 	428 
    -- CP-element group 419: successors 
    -- CP-element group 419: 	421 
    -- CP-element group 419:  members (3) 
      -- CP-element group 419: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_651_Update/cr
      -- CP-element group 419: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_651_Update/$entry
      -- CP-element group 419: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_651_update_start_
      -- 
    -- logger for CP element group try1_CP_1680_elements(419)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(419)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(419) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_651_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_4008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(419), ack => ADD_u12_u12_651_inst_req_1); -- 
    try1_cp_element_group_419: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_419"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(421) & try1_CP_1680_elements(440) & try1_CP_1680_elements(428);
      gj_try1_cp_element_group_419 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(419), clk => clk, reset => reset); --
    end block;
    -- CP-element group 420:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	418 
    -- CP-element group 420: successors 
    -- CP-element group 420: marked-successors 
    -- CP-element group 420: 	402 
    -- CP-element group 420: 	418 
    -- CP-element group 420:  members (3) 
      -- CP-element group 420: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_651_Sample/ra
      -- CP-element group 420: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_651_Sample/$exit
      -- CP-element group 420: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_651_sample_completed_
      -- 
    -- logger for CP element group try1_CP_1680_elements(420)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(420)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(420) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_651_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_651_inst_ack_0, ack => try1_CP_1680_elements(420)); -- 
    -- CP-element group 421:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	419 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	426 
    -- CP-element group 421: 	438 
    -- CP-element group 421: marked-successors 
    -- CP-element group 421: 	419 
    -- CP-element group 421:  members (29) 
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_651_Update/$exit
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_651_Update/ca
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_index_resize_0/index_resize_ack
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_index_scaled_0
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_index_resize_0/$exit
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_index_scale_0/$entry
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_word_address_calculated
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_index_scale_0/$exit
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_root_address_calculated
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_final_index_sum_regn/req
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_word_addrgen/root_register_req
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_word_addrgen/root_register_ack
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_offset_calculated
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_index_resized_0
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_final_index_sum_regn/$exit
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_word_addrgen/$exit
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_word_addrgen/$entry
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_651_update_completed_
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_base_plus_offset/sum_rename_ack
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_base_plus_offset/sum_rename_req
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_base_plus_offset/$exit
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_index_resize_0/$entry
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_base_plus_offset/$entry
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_index_resize_0/index_resize_req
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_final_index_sum_regn/ack
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_final_index_sum_regn/$entry
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_index_scale_0/scale_rename_ack
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_index_scale_0/scale_rename_req
      -- CP-element group 421: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_index_computed_0
      -- 
    -- logger for CP element group try1_CP_1680_elements(421)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(421)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(421) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_651_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_651_inst_ack_1, ack => try1_CP_1680_elements(421)); -- 
    -- CP-element group 422:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	404 
    -- CP-element group 422: marked-predecessors 
    -- CP-element group 422: 	424 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	424 
    -- CP-element group 422:  members (3) 
      -- CP-element group 422: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_655_sample_start_
      -- CP-element group 422: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_655_Sample/$entry
      -- CP-element group 422: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_655_Sample/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(422)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(422)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(422) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_H_574_delayed_5_0_653_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_4017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(422), ack => W_H_574_delayed_5_0_653_inst_req_0); -- 
    try1_cp_element_group_422: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_422"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(404) & try1_CP_1680_elements(424);
      gj_try1_cp_element_group_422 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(422), clk => clk, reset => reset); --
    end block;
    -- CP-element group 423:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: marked-predecessors 
    -- CP-element group 423: 	425 
    -- CP-element group 423: 	432 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	425 
    -- CP-element group 423:  members (3) 
      -- CP-element group 423: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_655_update_start_
      -- CP-element group 423: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_655_Update/$entry
      -- CP-element group 423: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_655_Update/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(423)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(423)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(423) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_H_574_delayed_5_0_653_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_4022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(423), ack => W_H_574_delayed_5_0_653_inst_req_1); -- 
    try1_cp_element_group_423: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_423"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(425) & try1_CP_1680_elements(432);
      gj_try1_cp_element_group_423 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(423), clk => clk, reset => reset); --
    end block;
    -- CP-element group 424:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	422 
    -- CP-element group 424: successors 
    -- CP-element group 424: marked-successors 
    -- CP-element group 424: 	402 
    -- CP-element group 424: 	422 
    -- CP-element group 424:  members (3) 
      -- CP-element group 424: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_655_sample_completed_
      -- CP-element group 424: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_655_Sample/$exit
      -- CP-element group 424: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_655_Sample/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(424)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(424)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(424) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_H_574_delayed_5_0_653_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_H_574_delayed_5_0_653_inst_ack_0, ack => try1_CP_1680_elements(424)); -- 
    -- CP-element group 425:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	423 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	430 
    -- CP-element group 425: marked-successors 
    -- CP-element group 425: 	423 
    -- CP-element group 425:  members (29) 
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_655_Update/ack
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_655_update_completed_
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_655_Update/$exit
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_word_address_calculated
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_root_address_calculated
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_offset_calculated
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_index_resized_0
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_index_scaled_0
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_index_computed_0
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_index_resize_0/$entry
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_index_resize_0/$exit
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_index_resize_0/index_resize_req
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_index_resize_0/index_resize_ack
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_index_scale_0/$entry
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_index_scale_0/$exit
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_index_scale_0/scale_rename_req
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_index_scale_0/scale_rename_ack
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_final_index_sum_regn/$entry
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_final_index_sum_regn/$exit
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_final_index_sum_regn/req
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_final_index_sum_regn/ack
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_base_plus_offset/$entry
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_base_plus_offset/$exit
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_base_plus_offset/sum_rename_req
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_base_plus_offset/sum_rename_ack
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_word_addrgen/$entry
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_word_addrgen/$exit
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_word_addrgen/root_register_req
      -- CP-element group 425: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(425)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(425)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(425) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_H_574_delayed_5_0_653_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_4023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 425_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_H_574_delayed_5_0_653_inst_ack_1, ack => try1_CP_1680_elements(425)); -- 
    -- CP-element group 426:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	421 
    -- CP-element group 426: marked-predecessors 
    -- CP-element group 426: 	464 
    -- CP-element group 426: 	428 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	428 
    -- CP-element group 426:  members (5) 
      -- CP-element group 426: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_Sample/word_access_start/word_0/rr
      -- CP-element group 426: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_Sample/word_access_start/$entry
      -- CP-element group 426: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_Sample/word_access_start/word_0/$entry
      -- CP-element group 426: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_sample_start_
      -- 
    -- logger for CP element group try1_CP_1680_elements(426)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(426)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(426) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_659_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(426), ack => array_obj_ref_659_load_0_req_0); -- 
    try1_cp_element_group_426: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_426"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(421) & try1_CP_1680_elements(464) & try1_CP_1680_elements(428);
      gj_try1_cp_element_group_426 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(426), clk => clk, reset => reset); --
    end block;
    -- CP-element group 427:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: marked-predecessors 
    -- CP-element group 427: 	429 
    -- CP-element group 427: 	432 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	429 
    -- CP-element group 427:  members (5) 
      -- CP-element group 427: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_update_start_
      -- CP-element group 427: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_Update/word_access_complete/word_0/$entry
      -- CP-element group 427: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_Update/$entry
      -- CP-element group 427: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_Update/word_access_complete/word_0/cr
      -- CP-element group 427: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_Update/word_access_complete/$entry
      -- 
    -- logger for CP element group try1_CP_1680_elements(427)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(427)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(427) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_659_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_4080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(427), ack => array_obj_ref_659_load_0_req_1); -- 
    try1_cp_element_group_427: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_427"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(429) & try1_CP_1680_elements(432);
      gj_try1_cp_element_group_427 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(427), clk => clk, reset => reset); --
    end block;
    -- CP-element group 428:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	426 
    -- CP-element group 428: successors 
    -- CP-element group 428: 	471 
    -- CP-element group 428: marked-successors 
    -- CP-element group 428: 	419 
    -- CP-element group 428: 	426 
    -- CP-element group 428:  members (5) 
      -- CP-element group 428: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_Sample/word_access_start/word_0/$exit
      -- CP-element group 428: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_Sample/word_access_start/$exit
      -- CP-element group 428: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_Sample/$exit
      -- CP-element group 428: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_sample_completed_
      -- CP-element group 428: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(428)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(428)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(428) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_659_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_659_load_0_ack_0, ack => try1_CP_1680_elements(428)); -- 
    -- CP-element group 429:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	427 
    -- CP-element group 429: successors 
    -- CP-element group 429: 	430 
    -- CP-element group 429: marked-successors 
    -- CP-element group 429: 	427 
    -- CP-element group 429:  members (9) 
      -- CP-element group 429: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_Update/word_access_complete/word_0/$exit
      -- CP-element group 429: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_Update/array_obj_ref_659_Merge/merge_req
      -- CP-element group 429: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_Update/array_obj_ref_659_Merge/merge_ack
      -- CP-element group 429: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_Update/$exit
      -- CP-element group 429: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_Update/word_access_complete/word_0/ca
      -- CP-element group 429: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_Update/array_obj_ref_659_Merge/$entry
      -- CP-element group 429: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_Update/array_obj_ref_659_Merge/$exit
      -- CP-element group 429: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_update_completed_
      -- CP-element group 429: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_Update/word_access_complete/$exit
      -- 
    -- logger for CP element group try1_CP_1680_elements(429)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(429)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(429) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_659_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 429_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_659_load_0_ack_1, ack => try1_CP_1680_elements(429)); -- 
    -- CP-element group 430:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	471 
    -- CP-element group 430: 	425 
    -- CP-element group 430: 	429 
    -- CP-element group 430: marked-predecessors 
    -- CP-element group 430: 	432 
    -- CP-element group 430: successors 
    -- CP-element group 430: 	432 
    -- CP-element group 430:  members (9) 
      -- CP-element group 430: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_sample_start_
      -- CP-element group 430: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_Sample/$entry
      -- CP-element group 430: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_Sample/array_obj_ref_657_Split/$entry
      -- CP-element group 430: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_Sample/array_obj_ref_657_Split/$exit
      -- CP-element group 430: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_Sample/array_obj_ref_657_Split/split_req
      -- CP-element group 430: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_Sample/array_obj_ref_657_Split/split_ack
      -- CP-element group 430: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_Sample/word_access_start/$entry
      -- CP-element group 430: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_Sample/word_access_start/word_0/$entry
      -- CP-element group 430: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(430)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(430)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(430) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_657_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(430), ack => array_obj_ref_657_store_0_req_0); -- 
    try1_cp_element_group_430: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_430"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= try1_CP_1680_elements(471) & try1_CP_1680_elements(425) & try1_CP_1680_elements(429) & try1_CP_1680_elements(432);
      gj_try1_cp_element_group_430 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(430), clk => clk, reset => reset); --
    end block;
    -- CP-element group 431:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: marked-predecessors 
    -- CP-element group 431: 	433 
    -- CP-element group 431: successors 
    -- CP-element group 431: 	433 
    -- CP-element group 431:  members (5) 
      -- CP-element group 431: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_update_start_
      -- CP-element group 431: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_Update/$entry
      -- CP-element group 431: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_Update/word_access_complete/$entry
      -- CP-element group 431: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_Update/word_access_complete/word_0/$entry
      -- CP-element group 431: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(431)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(431)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(431) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_657_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_4147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(431), ack => array_obj_ref_657_store_0_req_1); -- 
    try1_cp_element_group_431: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_431"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(433);
      gj_try1_cp_element_group_431 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(431), clk => clk, reset => reset); --
    end block;
    -- CP-element group 432:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	430 
    -- CP-element group 432: successors 
    -- CP-element group 432: 	472 
    -- CP-element group 432: marked-successors 
    -- CP-element group 432: 	423 
    -- CP-element group 432: 	427 
    -- CP-element group 432: 	430 
    -- CP-element group 432:  members (5) 
      -- CP-element group 432: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_sample_completed_
      -- CP-element group 432: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_Sample/$exit
      -- CP-element group 432: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_Sample/word_access_start/$exit
      -- CP-element group 432: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_Sample/word_access_start/word_0/$exit
      -- CP-element group 432: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(432)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(432)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(432) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_657_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_657_store_0_ack_0, ack => try1_CP_1680_elements(432)); -- 
    -- CP-element group 433:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	431 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	476 
    -- CP-element group 433: marked-successors 
    -- CP-element group 433: 	431 
    -- CP-element group 433:  members (5) 
      -- CP-element group 433: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_update_completed_
      -- CP-element group 433: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_Update/$exit
      -- CP-element group 433: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_Update/word_access_complete/$exit
      -- CP-element group 433: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_Update/word_access_complete/word_0/$exit
      -- CP-element group 433: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(433)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(433)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(433) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_657_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 433_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_657_store_0_ack_1, ack => try1_CP_1680_elements(433)); -- 
    -- CP-element group 434:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	404 
    -- CP-element group 434: marked-predecessors 
    -- CP-element group 434: 	436 
    -- CP-element group 434: successors 
    -- CP-element group 434: 	436 
    -- CP-element group 434:  members (3) 
      -- CP-element group 434: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_664_sample_start_
      -- CP-element group 434: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_664_Sample/$entry
      -- CP-element group 434: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_664_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(434)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(434)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(434) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_664_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(434), ack => ADD_u12_u12_664_inst_req_0); -- 
    try1_cp_element_group_434: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_434"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(404) & try1_CP_1680_elements(436);
      gj_try1_cp_element_group_434 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(434), clk => clk, reset => reset); --
    end block;
    -- CP-element group 435:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: marked-predecessors 
    -- CP-element group 435: 	456 
    -- CP-element group 435: 	444 
    -- CP-element group 435: 	437 
    -- CP-element group 435: successors 
    -- CP-element group 435: 	437 
    -- CP-element group 435:  members (3) 
      -- CP-element group 435: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_664_update_start_
      -- CP-element group 435: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_664_Update/$entry
      -- CP-element group 435: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_664_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(435)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(435)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(435) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_664_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_4161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(435), ack => ADD_u12_u12_664_inst_req_1); -- 
    try1_cp_element_group_435: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_435"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(456) & try1_CP_1680_elements(444) & try1_CP_1680_elements(437);
      gj_try1_cp_element_group_435 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(435), clk => clk, reset => reset); --
    end block;
    -- CP-element group 436:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	434 
    -- CP-element group 436: successors 
    -- CP-element group 436: marked-successors 
    -- CP-element group 436: 	402 
    -- CP-element group 436: 	434 
    -- CP-element group 436:  members (3) 
      -- CP-element group 436: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_664_sample_completed_
      -- CP-element group 436: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_664_Sample/$exit
      -- CP-element group 436: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_664_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(436)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(436)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(436) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_664_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 436_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_664_inst_ack_0, ack => try1_CP_1680_elements(436)); -- 
    -- CP-element group 437:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	435 
    -- CP-element group 437: successors 
    -- CP-element group 437: 	454 
    -- CP-element group 437: 	442 
    -- CP-element group 437: marked-successors 
    -- CP-element group 437: 	435 
    -- CP-element group 437:  members (29) 
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_664_update_completed_
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_664_Update/$exit
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_664_Update/ca
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_word_address_calculated
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_root_address_calculated
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_offset_calculated
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_index_resized_0
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_index_scaled_0
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_index_computed_0
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_index_resize_0/$entry
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_index_resize_0/$exit
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_index_resize_0/index_resize_req
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_index_resize_0/index_resize_ack
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_index_scale_0/$entry
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_index_scale_0/$exit
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_index_scale_0/scale_rename_req
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_index_scale_0/scale_rename_ack
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_final_index_sum_regn/$entry
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_final_index_sum_regn/$exit
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_final_index_sum_regn/req
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_final_index_sum_regn/ack
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_base_plus_offset/$entry
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_base_plus_offset/$exit
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_base_plus_offset/sum_rename_req
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_base_plus_offset/sum_rename_ack
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_word_addrgen/$entry
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_word_addrgen/$exit
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_word_addrgen/root_register_req
      -- CP-element group 437: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(437)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(437)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(437) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_664_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 437_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_664_inst_ack_1, ack => try1_CP_1680_elements(437)); -- 
    -- CP-element group 438:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	421 
    -- CP-element group 438: marked-predecessors 
    -- CP-element group 438: 	440 
    -- CP-element group 438: successors 
    -- CP-element group 438: 	440 
    -- CP-element group 438:  members (3) 
      -- CP-element group 438: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_668_sample_start_
      -- CP-element group 438: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_668_Sample/$entry
      -- CP-element group 438: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_668_Sample/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(438)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(438)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(438) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_HH_584_delayed_4_0_666_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_4170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(438), ack => W_HH_584_delayed_4_0_666_inst_req_0); -- 
    try1_cp_element_group_438: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_438"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(421) & try1_CP_1680_elements(440);
      gj_try1_cp_element_group_438 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(438), clk => clk, reset => reset); --
    end block;
    -- CP-element group 439:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: marked-predecessors 
    -- CP-element group 439: 	448 
    -- CP-element group 439: 	441 
    -- CP-element group 439: successors 
    -- CP-element group 439: 	441 
    -- CP-element group 439:  members (3) 
      -- CP-element group 439: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_668_update_start_
      -- CP-element group 439: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_668_Update/$entry
      -- CP-element group 439: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_668_Update/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(439)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(439)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(439) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_HH_584_delayed_4_0_666_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_4175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(439), ack => W_HH_584_delayed_4_0_666_inst_req_1); -- 
    try1_cp_element_group_439: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_439"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(448) & try1_CP_1680_elements(441);
      gj_try1_cp_element_group_439 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(439), clk => clk, reset => reset); --
    end block;
    -- CP-element group 440:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	438 
    -- CP-element group 440: successors 
    -- CP-element group 440: marked-successors 
    -- CP-element group 440: 	419 
    -- CP-element group 440: 	438 
    -- CP-element group 440:  members (3) 
      -- CP-element group 440: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_668_sample_completed_
      -- CP-element group 440: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_668_Sample/$exit
      -- CP-element group 440: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_668_Sample/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(440)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(440)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(440) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_HH_584_delayed_4_0_666_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 440_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_HH_584_delayed_4_0_666_inst_ack_0, ack => try1_CP_1680_elements(440)); -- 
    -- CP-element group 441:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	439 
    -- CP-element group 441: successors 
    -- CP-element group 441: 	446 
    -- CP-element group 441: marked-successors 
    -- CP-element group 441: 	439 
    -- CP-element group 441:  members (29) 
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_index_computed_0
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_668_update_completed_
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_668_Update/$exit
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_668_Update/ack
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_word_address_calculated
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_root_address_calculated
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_offset_calculated
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_index_resized_0
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_index_scaled_0
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_index_resize_0/$entry
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_index_resize_0/$exit
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_index_resize_0/index_resize_req
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_index_resize_0/index_resize_ack
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_index_scale_0/$entry
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_index_scale_0/$exit
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_index_scale_0/scale_rename_req
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_index_scale_0/scale_rename_ack
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_final_index_sum_regn/$entry
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_final_index_sum_regn/$exit
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_final_index_sum_regn/req
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_final_index_sum_regn/ack
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_base_plus_offset/$entry
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_base_plus_offset/$exit
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_base_plus_offset/sum_rename_req
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_base_plus_offset/sum_rename_ack
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_word_addrgen/$entry
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_word_addrgen/$exit
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_word_addrgen/root_register_req
      -- CP-element group 441: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(441)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(441)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(441) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_HH_584_delayed_4_0_666_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_4176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 441_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_HH_584_delayed_4_0_666_inst_ack_1, ack => try1_CP_1680_elements(441)); -- 
    -- CP-element group 442:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	472 
    -- CP-element group 442: 	437 
    -- CP-element group 442: marked-predecessors 
    -- CP-element group 442: 	444 
    -- CP-element group 442: successors 
    -- CP-element group 442: 	444 
    -- CP-element group 442:  members (5) 
      -- CP-element group 442: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_sample_start_
      -- CP-element group 442: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_Sample/$entry
      -- CP-element group 442: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_Sample/word_access_start/$entry
      -- CP-element group 442: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_Sample/word_access_start/word_0/$entry
      -- CP-element group 442: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(442)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(442)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(442) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_672_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(442), ack => array_obj_ref_672_load_0_req_0); -- 
    try1_cp_element_group_442: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_442"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(472) & try1_CP_1680_elements(437) & try1_CP_1680_elements(444);
      gj_try1_cp_element_group_442 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(442), clk => clk, reset => reset); --
    end block;
    -- CP-element group 443:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: marked-predecessors 
    -- CP-element group 443: 	448 
    -- CP-element group 443: 	445 
    -- CP-element group 443: successors 
    -- CP-element group 443: 	445 
    -- CP-element group 443:  members (5) 
      -- CP-element group 443: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_update_start_
      -- CP-element group 443: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_Update/$entry
      -- CP-element group 443: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_Update/word_access_complete/$entry
      -- CP-element group 443: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_Update/word_access_complete/word_0/$entry
      -- CP-element group 443: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(443)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(443)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(443) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_672_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_4233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(443), ack => array_obj_ref_672_load_0_req_1); -- 
    try1_cp_element_group_443: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_443"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(448) & try1_CP_1680_elements(445);
      gj_try1_cp_element_group_443 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(443), clk => clk, reset => reset); --
    end block;
    -- CP-element group 444:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	442 
    -- CP-element group 444: successors 
    -- CP-element group 444: 	473 
    -- CP-element group 444: marked-successors 
    -- CP-element group 444: 	442 
    -- CP-element group 444: 	435 
    -- CP-element group 444:  members (5) 
      -- CP-element group 444: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_sample_completed_
      -- CP-element group 444: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_Sample/$exit
      -- CP-element group 444: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_Sample/word_access_start/$exit
      -- CP-element group 444: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_Sample/word_access_start/word_0/$exit
      -- CP-element group 444: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(444)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(444)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(444) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_672_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 444_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_672_load_0_ack_0, ack => try1_CP_1680_elements(444)); -- 
    -- CP-element group 445:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	443 
    -- CP-element group 445: successors 
    -- CP-element group 445: 	446 
    -- CP-element group 445: marked-successors 
    -- CP-element group 445: 	443 
    -- CP-element group 445:  members (9) 
      -- CP-element group 445: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_update_completed_
      -- CP-element group 445: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_Update/$exit
      -- CP-element group 445: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_Update/word_access_complete/$exit
      -- CP-element group 445: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_Update/word_access_complete/word_0/$exit
      -- CP-element group 445: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_Update/word_access_complete/word_0/ca
      -- CP-element group 445: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_Update/array_obj_ref_672_Merge/$entry
      -- CP-element group 445: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_Update/array_obj_ref_672_Merge/$exit
      -- CP-element group 445: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_Update/array_obj_ref_672_Merge/merge_req
      -- CP-element group 445: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_Update/array_obj_ref_672_Merge/merge_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(445)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(445)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(445) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_672_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 445_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_672_load_0_ack_1, ack => try1_CP_1680_elements(445)); -- 
    -- CP-element group 446:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	473 
    -- CP-element group 446: 	441 
    -- CP-element group 446: 	445 
    -- CP-element group 446: marked-predecessors 
    -- CP-element group 446: 	448 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	448 
    -- CP-element group 446:  members (9) 
      -- CP-element group 446: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_sample_start_
      -- CP-element group 446: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_Sample/$entry
      -- CP-element group 446: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_Sample/array_obj_ref_670_Split/$entry
      -- CP-element group 446: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_Sample/array_obj_ref_670_Split/$exit
      -- CP-element group 446: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_Sample/array_obj_ref_670_Split/split_req
      -- CP-element group 446: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_Sample/array_obj_ref_670_Split/split_ack
      -- CP-element group 446: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_Sample/word_access_start/$entry
      -- CP-element group 446: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_Sample/word_access_start/word_0/$entry
      -- CP-element group 446: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(446)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(446)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(446) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_670_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(446), ack => array_obj_ref_670_store_0_req_0); -- 
    try1_cp_element_group_446: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_446"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= try1_CP_1680_elements(473) & try1_CP_1680_elements(441) & try1_CP_1680_elements(445) & try1_CP_1680_elements(448);
      gj_try1_cp_element_group_446 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(446), clk => clk, reset => reset); --
    end block;
    -- CP-element group 447:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: marked-predecessors 
    -- CP-element group 447: 	449 
    -- CP-element group 447: successors 
    -- CP-element group 447: 	449 
    -- CP-element group 447:  members (5) 
      -- CP-element group 447: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_update_start_
      -- CP-element group 447: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_Update/$entry
      -- CP-element group 447: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_Update/word_access_complete/$entry
      -- CP-element group 447: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_Update/word_access_complete/word_0/$entry
      -- CP-element group 447: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(447)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(447)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(447) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_670_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_4300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(447), ack => array_obj_ref_670_store_0_req_1); -- 
    try1_cp_element_group_447: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_447"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(449);
      gj_try1_cp_element_group_447 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(447), clk => clk, reset => reset); --
    end block;
    -- CP-element group 448:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	446 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	474 
    -- CP-element group 448: marked-successors 
    -- CP-element group 448: 	443 
    -- CP-element group 448: 	439 
    -- CP-element group 448: 	446 
    -- CP-element group 448:  members (5) 
      -- CP-element group 448: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_sample_completed_
      -- CP-element group 448: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_Sample/$exit
      -- CP-element group 448: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_Sample/word_access_start/$exit
      -- CP-element group 448: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_Sample/word_access_start/word_0/$exit
      -- CP-element group 448: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(448)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(448)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(448) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_670_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 448_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_670_store_0_ack_0, ack => try1_CP_1680_elements(448)); -- 
    -- CP-element group 449:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	447 
    -- CP-element group 449: successors 
    -- CP-element group 449: 	476 
    -- CP-element group 449: marked-successors 
    -- CP-element group 449: 	447 
    -- CP-element group 449:  members (5) 
      -- CP-element group 449: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_update_completed_
      -- CP-element group 449: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_Update/$exit
      -- CP-element group 449: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_Update/word_access_complete/$exit
      -- CP-element group 449: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_Update/word_access_complete/word_0/$exit
      -- CP-element group 449: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(449)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(449)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(449) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_670_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 449_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_670_store_0_ack_1, ack => try1_CP_1680_elements(449)); -- 
    -- CP-element group 450:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	404 
    -- CP-element group 450: marked-predecessors 
    -- CP-element group 450: 	452 
    -- CP-element group 450: successors 
    -- CP-element group 450: 	452 
    -- CP-element group 450:  members (3) 
      -- CP-element group 450: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_677_sample_start_
      -- CP-element group 450: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_677_Sample/$entry
      -- CP-element group 450: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_677_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(450)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(450)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(450) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_677_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(450), ack => ADD_u12_u12_677_inst_req_0); -- 
    try1_cp_element_group_450: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_450"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(404) & try1_CP_1680_elements(452);
      gj_try1_cp_element_group_450 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(450), clk => clk, reset => reset); --
    end block;
    -- CP-element group 451:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: marked-predecessors 
    -- CP-element group 451: 	460 
    -- CP-element group 451: 	453 
    -- CP-element group 451: successors 
    -- CP-element group 451: 	453 
    -- CP-element group 451:  members (3) 
      -- CP-element group 451: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_677_update_start_
      -- CP-element group 451: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_677_Update/$entry
      -- CP-element group 451: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_677_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(451)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(451)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(451) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_677_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_4314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(451), ack => ADD_u12_u12_677_inst_req_1); -- 
    try1_cp_element_group_451: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_451"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(460) & try1_CP_1680_elements(453);
      gj_try1_cp_element_group_451 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(451), clk => clk, reset => reset); --
    end block;
    -- CP-element group 452:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	450 
    -- CP-element group 452: successors 
    -- CP-element group 452: marked-successors 
    -- CP-element group 452: 	450 
    -- CP-element group 452: 	402 
    -- CP-element group 452:  members (3) 
      -- CP-element group 452: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_677_sample_completed_
      -- CP-element group 452: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_677_Sample/$exit
      -- CP-element group 452: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_677_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(452)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(452)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(452) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_677_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 452_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_677_inst_ack_0, ack => try1_CP_1680_elements(452)); -- 
    -- CP-element group 453:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	451 
    -- CP-element group 453: successors 
    -- CP-element group 453: 	458 
    -- CP-element group 453: marked-successors 
    -- CP-element group 453: 	451 
    -- CP-element group 453:  members (29) 
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_677_update_completed_
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_677_Update/$exit
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_677_Update/ca
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_word_address_calculated
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_root_address_calculated
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_offset_calculated
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_index_resized_0
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_index_scaled_0
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_index_computed_0
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_index_resize_0/$entry
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_index_resize_0/$exit
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_index_resize_0/index_resize_req
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_index_resize_0/index_resize_ack
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_index_scale_0/$entry
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_index_scale_0/$exit
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_index_scale_0/scale_rename_req
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_index_scale_0/scale_rename_ack
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_final_index_sum_regn/$entry
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_final_index_sum_regn/$exit
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_final_index_sum_regn/req
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_final_index_sum_regn/ack
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_base_plus_offset/$entry
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_base_plus_offset/$exit
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_base_plus_offset/sum_rename_req
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_base_plus_offset/sum_rename_ack
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_word_addrgen/$entry
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_word_addrgen/$exit
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_word_addrgen/root_register_req
      -- CP-element group 453: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(453)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(453)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(453) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_677_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 453_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_677_inst_ack_1, ack => try1_CP_1680_elements(453)); -- 
    -- CP-element group 454:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	437 
    -- CP-element group 454: marked-predecessors 
    -- CP-element group 454: 	456 
    -- CP-element group 454: successors 
    -- CP-element group 454: 	456 
    -- CP-element group 454:  members (3) 
      -- CP-element group 454: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_681_sample_start_
      -- CP-element group 454: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_681_Sample/$entry
      -- CP-element group 454: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_681_Sample/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(454)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(454)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(454) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_HHH_594_delayed_4_0_679_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_4323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(454), ack => W_HHH_594_delayed_4_0_679_inst_req_0); -- 
    try1_cp_element_group_454: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_454"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(437) & try1_CP_1680_elements(456);
      gj_try1_cp_element_group_454 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(454), clk => clk, reset => reset); --
    end block;
    -- CP-element group 455:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: marked-predecessors 
    -- CP-element group 455: 	457 
    -- CP-element group 455: 	464 
    -- CP-element group 455: successors 
    -- CP-element group 455: 	457 
    -- CP-element group 455:  members (3) 
      -- CP-element group 455: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_681_update_start_
      -- CP-element group 455: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_681_Update/$entry
      -- CP-element group 455: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_681_Update/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(455)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(455)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(455) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_HHH_594_delayed_4_0_679_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_4328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(455), ack => W_HHH_594_delayed_4_0_679_inst_req_1); -- 
    try1_cp_element_group_455: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_455"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(457) & try1_CP_1680_elements(464);
      gj_try1_cp_element_group_455 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(455), clk => clk, reset => reset); --
    end block;
    -- CP-element group 456:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	454 
    -- CP-element group 456: successors 
    -- CP-element group 456: marked-successors 
    -- CP-element group 456: 	454 
    -- CP-element group 456: 	435 
    -- CP-element group 456:  members (3) 
      -- CP-element group 456: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_681_sample_completed_
      -- CP-element group 456: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_681_Sample/$exit
      -- CP-element group 456: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_681_Sample/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(456)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(456)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(456) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_HHH_594_delayed_4_0_679_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 456_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_HHH_594_delayed_4_0_679_inst_ack_0, ack => try1_CP_1680_elements(456)); -- 
    -- CP-element group 457:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	455 
    -- CP-element group 457: successors 
    -- CP-element group 457: 	462 
    -- CP-element group 457: marked-successors 
    -- CP-element group 457: 	455 
    -- CP-element group 457:  members (29) 
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_681_update_completed_
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_681_Update/$exit
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/assign_stmt_681_Update/ack
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_word_address_calculated
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_root_address_calculated
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_offset_calculated
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_index_resized_0
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_index_scaled_0
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_index_computed_0
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_index_resize_0/$entry
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_index_resize_0/$exit
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_index_resize_0/index_resize_req
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_index_resize_0/index_resize_ack
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_index_scale_0/$entry
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_index_scale_0/$exit
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_index_scale_0/scale_rename_req
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_index_scale_0/scale_rename_ack
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_final_index_sum_regn/$entry
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_final_index_sum_regn/$exit
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_final_index_sum_regn/req
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_final_index_sum_regn/ack
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_base_plus_offset/$entry
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_base_plus_offset/$exit
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_base_plus_offset/sum_rename_req
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_base_plus_offset/sum_rename_ack
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_word_addrgen/$entry
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_word_addrgen/$exit
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_word_addrgen/root_register_req
      -- CP-element group 457: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(457)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(457)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(457) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:W_HHH_594_delayed_4_0_679_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_4329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 457_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_HHH_594_delayed_4_0_679_inst_ack_1, ack => try1_CP_1680_elements(457)); -- 
    -- CP-element group 458:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	474 
    -- CP-element group 458: 	453 
    -- CP-element group 458: marked-predecessors 
    -- CP-element group 458: 	460 
    -- CP-element group 458: successors 
    -- CP-element group 458: 	460 
    -- CP-element group 458:  members (5) 
      -- CP-element group 458: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_sample_start_
      -- CP-element group 458: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_Sample/$entry
      -- CP-element group 458: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_Sample/word_access_start/$entry
      -- CP-element group 458: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_Sample/word_access_start/word_0/$entry
      -- CP-element group 458: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(458)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(458)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(458) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_685_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(458), ack => array_obj_ref_685_load_0_req_0); -- 
    try1_cp_element_group_458: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_458"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(474) & try1_CP_1680_elements(453) & try1_CP_1680_elements(460);
      gj_try1_cp_element_group_458 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(458), clk => clk, reset => reset); --
    end block;
    -- CP-element group 459:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: marked-predecessors 
    -- CP-element group 459: 	461 
    -- CP-element group 459: 	464 
    -- CP-element group 459: successors 
    -- CP-element group 459: 	461 
    -- CP-element group 459:  members (5) 
      -- CP-element group 459: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_update_start_
      -- CP-element group 459: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_Update/$entry
      -- CP-element group 459: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_Update/word_access_complete/$entry
      -- CP-element group 459: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_Update/word_access_complete/word_0/$entry
      -- CP-element group 459: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(459)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(459)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(459) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_685_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_4386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(459), ack => array_obj_ref_685_load_0_req_1); -- 
    try1_cp_element_group_459: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_459"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(461) & try1_CP_1680_elements(464);
      gj_try1_cp_element_group_459 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(459), clk => clk, reset => reset); --
    end block;
    -- CP-element group 460:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: 	458 
    -- CP-element group 460: successors 
    -- CP-element group 460: 	475 
    -- CP-element group 460: marked-successors 
    -- CP-element group 460: 	458 
    -- CP-element group 460: 	451 
    -- CP-element group 460:  members (5) 
      -- CP-element group 460: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_sample_completed_
      -- CP-element group 460: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_Sample/$exit
      -- CP-element group 460: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_Sample/word_access_start/$exit
      -- CP-element group 460: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_Sample/word_access_start/word_0/$exit
      -- CP-element group 460: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(460)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(460)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(460) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_685_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 460_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_685_load_0_ack_0, ack => try1_CP_1680_elements(460)); -- 
    -- CP-element group 461:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: 	459 
    -- CP-element group 461: successors 
    -- CP-element group 461: 	462 
    -- CP-element group 461: marked-successors 
    -- CP-element group 461: 	459 
    -- CP-element group 461:  members (9) 
      -- CP-element group 461: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_update_completed_
      -- CP-element group 461: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_Update/$exit
      -- CP-element group 461: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_Update/word_access_complete/$exit
      -- CP-element group 461: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_Update/word_access_complete/word_0/$exit
      -- CP-element group 461: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_Update/word_access_complete/word_0/ca
      -- CP-element group 461: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_Update/array_obj_ref_685_Merge/$entry
      -- CP-element group 461: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_Update/array_obj_ref_685_Merge/$exit
      -- CP-element group 461: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_Update/array_obj_ref_685_Merge/merge_req
      -- CP-element group 461: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_Update/array_obj_ref_685_Merge/merge_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(461)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(461)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(461) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_685_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 461_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_685_load_0_ack_1, ack => try1_CP_1680_elements(461)); -- 
    -- CP-element group 462:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: 	475 
    -- CP-element group 462: 	461 
    -- CP-element group 462: 	457 
    -- CP-element group 462: marked-predecessors 
    -- CP-element group 462: 	464 
    -- CP-element group 462: successors 
    -- CP-element group 462: 	464 
    -- CP-element group 462:  members (9) 
      -- CP-element group 462: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_sample_start_
      -- CP-element group 462: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_Sample/$entry
      -- CP-element group 462: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_Sample/array_obj_ref_683_Split/$entry
      -- CP-element group 462: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_Sample/array_obj_ref_683_Split/$exit
      -- CP-element group 462: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_Sample/array_obj_ref_683_Split/split_req
      -- CP-element group 462: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_Sample/array_obj_ref_683_Split/split_ack
      -- CP-element group 462: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_Sample/word_access_start/$entry
      -- CP-element group 462: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_Sample/word_access_start/word_0/$entry
      -- CP-element group 462: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(462)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(462)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(462) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_683_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(462), ack => array_obj_ref_683_store_0_req_0); -- 
    try1_cp_element_group_462: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_462"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= try1_CP_1680_elements(475) & try1_CP_1680_elements(461) & try1_CP_1680_elements(457) & try1_CP_1680_elements(464);
      gj_try1_cp_element_group_462 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(462), clk => clk, reset => reset); --
    end block;
    -- CP-element group 463:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: marked-predecessors 
    -- CP-element group 463: 	465 
    -- CP-element group 463: successors 
    -- CP-element group 463: 	465 
    -- CP-element group 463:  members (5) 
      -- CP-element group 463: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_update_start_
      -- CP-element group 463: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_Update/$entry
      -- CP-element group 463: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_Update/word_access_complete/$entry
      -- CP-element group 463: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_Update/word_access_complete/word_0/$entry
      -- CP-element group 463: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(463)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(463)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(463) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_683_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_4453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(463), ack => array_obj_ref_683_store_0_req_1); -- 
    try1_cp_element_group_463: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_463"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= try1_CP_1680_elements(465);
      gj_try1_cp_element_group_463 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(463), clk => clk, reset => reset); --
    end block;
    -- CP-element group 464:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: 	462 
    -- CP-element group 464: successors 
    -- CP-element group 464: 	476 
    -- CP-element group 464: marked-successors 
    -- CP-element group 464: 	462 
    -- CP-element group 464: 	459 
    -- CP-element group 464: 	455 
    -- CP-element group 464: 	426 
    -- CP-element group 464:  members (6) 
      -- CP-element group 464: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_sample_completed_
      -- CP-element group 464: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_Sample/$exit
      -- CP-element group 464: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_Sample/word_access_start/$exit
      -- CP-element group 464: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_Sample/word_access_start/word_0/$exit
      -- CP-element group 464: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_Sample/word_access_start/word_0/ra
      -- CP-element group 464: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ring_reenable_memory_space_3
      -- 
    -- logger for CP element group try1_CP_1680_elements(464)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(464)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(464) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_683_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 464_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_683_store_0_ack_0, ack => try1_CP_1680_elements(464)); -- 
    -- CP-element group 465:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: 	463 
    -- CP-element group 465: successors 
    -- CP-element group 465: 	476 
    -- CP-element group 465: marked-successors 
    -- CP-element group 465: 	463 
    -- CP-element group 465:  members (5) 
      -- CP-element group 465: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_update_completed_
      -- CP-element group 465: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_Update/$exit
      -- CP-element group 465: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_Update/word_access_complete/$exit
      -- CP-element group 465: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_Update/word_access_complete/word_0/$exit
      -- CP-element group 465: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_683_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(465)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(465)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(465) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_683_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 465_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_683_store_0_ack_1, ack => try1_CP_1680_elements(465)); -- 
    -- CP-element group 466:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: 	404 
    -- CP-element group 466: marked-predecessors 
    -- CP-element group 466: 	468 
    -- CP-element group 466: successors 
    -- CP-element group 466: 	468 
    -- CP-element group 466:  members (3) 
      -- CP-element group 466: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_690_sample_start_
      -- CP-element group 466: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_690_Sample/$entry
      -- CP-element group 466: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_690_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(466)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(466)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(466) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_690_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(466), ack => ADD_u12_u12_690_inst_req_0); -- 
    try1_cp_element_group_466: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 25) := "try1_cp_element_group_466"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(404) & try1_CP_1680_elements(468);
      gj_try1_cp_element_group_466 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(466), clk => clk, reset => reset); --
    end block;
    -- CP-element group 467:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: 	403 
    -- CP-element group 467: marked-predecessors 
    -- CP-element group 467: 	469 
    -- CP-element group 467: successors 
    -- CP-element group 467: 	469 
    -- CP-element group 467:  members (3) 
      -- CP-element group 467: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_690_update_start_
      -- CP-element group 467: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_690_Update/$entry
      -- CP-element group 467: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_690_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(467)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(467)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(467) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_690_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_4467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(467), ack => ADD_u12_u12_690_inst_req_1); -- 
    try1_cp_element_group_467: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_467"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(403) & try1_CP_1680_elements(469);
      gj_try1_cp_element_group_467 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(467), clk => clk, reset => reset); --
    end block;
    -- CP-element group 468:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: 	466 
    -- CP-element group 468: successors 
    -- CP-element group 468: marked-successors 
    -- CP-element group 468: 	402 
    -- CP-element group 468: 	466 
    -- CP-element group 468:  members (3) 
      -- CP-element group 468: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_690_sample_completed_
      -- CP-element group 468: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_690_Sample/$exit
      -- CP-element group 468: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_690_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(468)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(468)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(468) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_690_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 468_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_690_inst_ack_0, ack => try1_CP_1680_elements(468)); -- 
    -- CP-element group 469:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: 	467 
    -- CP-element group 469: successors 
    -- CP-element group 469: 	399 
    -- CP-element group 469: marked-successors 
    -- CP-element group 469: 	401 
    -- CP-element group 469: 	467 
    -- CP-element group 469:  members (3) 
      -- CP-element group 469: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_690_update_completed_
      -- CP-element group 469: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_690_Update/$exit
      -- CP-element group 469: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/ADD_u12_u12_690_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(469)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(469)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(469) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_690_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 469_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_690_inst_ack_1, ack => try1_CP_1680_elements(469)); -- 
    -- CP-element group 470:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: 	398 
    -- CP-element group 470: successors 
    -- CP-element group 470: 	399 
    -- CP-element group 470:  members (1) 
      -- CP-element group 470: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group try1_CP_1680_elements(470)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(470)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(470) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(470) is a control-delay.
    cp_element_470_delay: control_delay_element  generic map(name => " 470_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(398), ack => try1_CP_1680_elements(470), clk => clk, reset =>reset);
    -- CP-element group 471:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: 	428 
    -- CP-element group 471: successors 
    -- CP-element group 471: 	430 
    -- CP-element group 471:  members (1) 
      -- CP-element group 471: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_659_array_obj_ref_657_delay
      -- 
    -- logger for CP element group try1_CP_1680_elements(471)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(471)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(471) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(471) is a control-delay.
    cp_element_471_delay: control_delay_element  generic map(name => " 471_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(428), ack => try1_CP_1680_elements(471), clk => clk, reset =>reset);
    -- CP-element group 472:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: 	432 
    -- CP-element group 472: successors 
    -- CP-element group 472: 	442 
    -- CP-element group 472:  members (1) 
      -- CP-element group 472: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_657_array_obj_ref_672_delay
      -- 
    -- logger for CP element group try1_CP_1680_elements(472)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(472)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(472) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(472) is a control-delay.
    cp_element_472_delay: control_delay_element  generic map(name => " 472_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(432), ack => try1_CP_1680_elements(472), clk => clk, reset =>reset);
    -- CP-element group 473:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	444 
    -- CP-element group 473: successors 
    -- CP-element group 473: 	446 
    -- CP-element group 473:  members (1) 
      -- CP-element group 473: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_672_array_obj_ref_670_delay
      -- 
    -- logger for CP element group try1_CP_1680_elements(473)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(473)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(473) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(473) is a control-delay.
    cp_element_473_delay: control_delay_element  generic map(name => " 473_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(444), ack => try1_CP_1680_elements(473), clk => clk, reset =>reset);
    -- CP-element group 474:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	448 
    -- CP-element group 474: successors 
    -- CP-element group 474: 	458 
    -- CP-element group 474:  members (1) 
      -- CP-element group 474: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_670_array_obj_ref_685_delay
      -- 
    -- logger for CP element group try1_CP_1680_elements(474)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(474)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(474) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(474) is a control-delay.
    cp_element_474_delay: control_delay_element  generic map(name => " 474_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(448), ack => try1_CP_1680_elements(474), clk => clk, reset =>reset);
    -- CP-element group 475:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: 	460 
    -- CP-element group 475: successors 
    -- CP-element group 475: 	462 
    -- CP-element group 475:  members (1) 
      -- CP-element group 475: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/array_obj_ref_685_array_obj_ref_683_delay
      -- 
    -- logger for CP element group try1_CP_1680_elements(475)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(475)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(475) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(475) is a control-delay.
    cp_element_475_delay: control_delay_element  generic map(name => " 475_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(460), ack => try1_CP_1680_elements(475), clk => clk, reset =>reset);
    -- CP-element group 476:  join  transition  bypass  pipeline-parent 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: 	449 
    -- CP-element group 476: 	433 
    -- CP-element group 476: 	464 
    -- CP-element group 476: 	465 
    -- CP-element group 476: successors 
    -- CP-element group 476: 	395 
    -- CP-element group 476:  members (1) 
      -- CP-element group 476: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/do_while_stmt_640_loop_body/$exit
      -- 
    -- logger for CP element group try1_CP_1680_elements(476)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(476)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(476) fired."); 
        -- 
      end if; --
    end process; 
    try1_cp_element_group_476: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 7,2 => 7,3 => 7);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_476"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= try1_CP_1680_elements(449) & try1_CP_1680_elements(433) & try1_CP_1680_elements(464) & try1_CP_1680_elements(465);
      gj_try1_cp_element_group_476 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(476), clk => clk, reset => reset); --
    end block;
    -- CP-element group 477:  transition  input  bypass  pipeline-parent 
    -- CP-element group 477: predecessors 
    -- CP-element group 477: 	394 
    -- CP-element group 477: successors 
    -- CP-element group 477:  members (2) 
      -- CP-element group 477: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/loop_exit/$exit
      -- CP-element group 477: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/loop_exit/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(477)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(477)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(477) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:do_while_stmt_640_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 477_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_640_branch_ack_0, ack => try1_CP_1680_elements(477)); -- 
    -- CP-element group 478:  transition  input  bypass  pipeline-parent 
    -- CP-element group 478: predecessors 
    -- CP-element group 478: 	394 
    -- CP-element group 478: successors 
    -- CP-element group 478:  members (2) 
      -- CP-element group 478: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/loop_taken/$exit
      -- CP-element group 478: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/loop_taken/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(478)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(478)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(478) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:do_while_stmt_640_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_4483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 478_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_640_branch_ack_1, ack => try1_CP_1680_elements(478)); -- 
    -- CP-element group 479:  transition  bypass  pipeline-parent 
    -- CP-element group 479: predecessors 
    -- CP-element group 479: 	392 
    -- CP-element group 479: successors 
    -- CP-element group 479: 	390 
    -- CP-element group 479:  members (1) 
      -- CP-element group 479: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_639/do_while_stmt_640/$exit
      -- 
    -- logger for CP element group try1_CP_1680_elements(479)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(479)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(479) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(479) <= try1_CP_1680_elements(392);
    -- CP-element group 480:  transition  input  bypass 
    -- CP-element group 480: predecessors 
    -- CP-element group 480: 	390 
    -- CP-element group 480: successors 
    -- CP-element group 480:  members (3) 
      -- CP-element group 480: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_702_sample_completed_
      -- CP-element group 480: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_702_Sample/$exit
      -- CP-element group 480: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_702_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(480)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(480)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(480) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_702_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 480_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_702_inst_ack_0, ack => try1_CP_1680_elements(480)); -- 
    -- CP-element group 481:  transition  input  output  bypass 
    -- CP-element group 481: predecessors 
    -- CP-element group 481: 	390 
    -- CP-element group 481: successors 
    -- CP-element group 481: 	482 
    -- CP-element group 481:  members (6) 
      -- CP-element group 481: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/call_stmt_705_sample_start_
      -- CP-element group 481: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_702_update_completed_
      -- CP-element group 481: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_702_Update/$exit
      -- CP-element group 481: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_702_Update/ca
      -- CP-element group 481: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/call_stmt_705_Sample/$entry
      -- CP-element group 481: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/call_stmt_705_Sample/crr
      -- 
    -- logger for CP element group try1_CP_1680_elements(481)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(481)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(481) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_702_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:call_stmt_705_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_4505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 481_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_702_inst_ack_1, ack => try1_CP_1680_elements(481)); -- 
    crr_4509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(481), ack => call_stmt_705_call_req_0); -- 
    -- CP-element group 482:  transition  input  bypass 
    -- CP-element group 482: predecessors 
    -- CP-element group 482: 	481 
    -- CP-element group 482: successors 
    -- CP-element group 482:  members (3) 
      -- CP-element group 482: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/call_stmt_705_sample_completed_
      -- CP-element group 482: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/call_stmt_705_Sample/$exit
      -- CP-element group 482: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/call_stmt_705_Sample/cra
      -- 
    -- logger for CP element group try1_CP_1680_elements(482)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(482)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(482) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:call_stmt_705_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_4510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 482_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_705_call_ack_0, ack => try1_CP_1680_elements(482)); -- 
    -- CP-element group 483:  fork  transition  input  output  bypass 
    -- CP-element group 483: predecessors 
    -- CP-element group 483: 	390 
    -- CP-element group 483: successors 
    -- CP-element group 483: 	484 
    -- CP-element group 483: 	494 
    -- CP-element group 483: 	499 
    -- CP-element group 483: 	489 
    -- CP-element group 483:  members (15) 
      -- CP-element group 483: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/call_stmt_705_update_completed_
      -- CP-element group 483: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/call_stmt_705_Update/$exit
      -- CP-element group 483: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/call_stmt_705_Update/cca
      -- CP-element group 483: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_709_sample_start_
      -- CP-element group 483: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_709_Sample/$entry
      -- CP-element group 483: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_709_Sample/rr
      -- CP-element group 483: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_714_sample_start_
      -- CP-element group 483: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_714_Sample/$entry
      -- CP-element group 483: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_714_Sample/rr
      -- CP-element group 483: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_719_sample_start_
      -- CP-element group 483: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_719_Sample/$entry
      -- CP-element group 483: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_719_Sample/rr
      -- CP-element group 483: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_724_sample_start_
      -- CP-element group 483: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_724_Sample/$entry
      -- CP-element group 483: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_724_Sample/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(483)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(483)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(483) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:call_stmt_705_call_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_709_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_719_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_724_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_714_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    cca_4515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 483_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_705_call_ack_1, ack => try1_CP_1680_elements(483)); -- 
    rr_4523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(483), ack => slice_709_inst_req_0); -- 
    rr_4617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(483), ack => slice_719_inst_req_0); -- 
    rr_4664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(483), ack => slice_724_inst_req_0); -- 
    rr_4570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(483), ack => slice_714_inst_req_0); -- 
    -- CP-element group 484:  transition  input  bypass 
    -- CP-element group 484: predecessors 
    -- CP-element group 484: 	483 
    -- CP-element group 484: successors 
    -- CP-element group 484:  members (3) 
      -- CP-element group 484: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_709_sample_completed_
      -- CP-element group 484: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_709_Sample/$exit
      -- CP-element group 484: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_709_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(484)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(484)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(484) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_709_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 484_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_709_inst_ack_0, ack => try1_CP_1680_elements(484)); -- 
    -- CP-element group 485:  transition  input  bypass 
    -- CP-element group 485: predecessors 
    -- CP-element group 485: 	390 
    -- CP-element group 485: successors 
    -- CP-element group 485: 	486 
    -- CP-element group 485:  members (3) 
      -- CP-element group 485: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_709_update_completed_
      -- CP-element group 485: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_709_Update/$exit
      -- CP-element group 485: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_709_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(485)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(485)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(485) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_709_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 485_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_709_inst_ack_1, ack => try1_CP_1680_elements(485)); -- 
    -- CP-element group 486:  join  transition  output  bypass 
    -- CP-element group 486: predecessors 
    -- CP-element group 486: 	485 
    -- CP-element group 486: 	390 
    -- CP-element group 486: successors 
    -- CP-element group 486: 	487 
    -- CP-element group 486:  members (9) 
      -- CP-element group 486: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_sample_start_
      -- CP-element group 486: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_Sample/$entry
      -- CP-element group 486: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_Sample/array_obj_ref_707_Split/$entry
      -- CP-element group 486: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_Sample/array_obj_ref_707_Split/$exit
      -- CP-element group 486: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_Sample/array_obj_ref_707_Split/split_req
      -- CP-element group 486: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_Sample/array_obj_ref_707_Split/split_ack
      -- CP-element group 486: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_Sample/word_access_start/$entry
      -- CP-element group 486: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_Sample/word_access_start/word_0/$entry
      -- CP-element group 486: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(486)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(486)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(486) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_707_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(486), ack => array_obj_ref_707_store_0_req_0); -- 
    try1_cp_element_group_486: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_486"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(485) & try1_CP_1680_elements(390);
      gj_try1_cp_element_group_486 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(486), clk => clk, reset => reset); --
    end block;
    -- CP-element group 487:  transition  input  bypass 
    -- CP-element group 487: predecessors 
    -- CP-element group 487: 	486 
    -- CP-element group 487: successors 
    -- CP-element group 487: 	506 
    -- CP-element group 487:  members (5) 
      -- CP-element group 487: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_sample_completed_
      -- CP-element group 487: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_Sample/$exit
      -- CP-element group 487: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_Sample/word_access_start/$exit
      -- CP-element group 487: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_Sample/word_access_start/word_0/$exit
      -- CP-element group 487: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(487)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(487)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(487) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_707_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 487_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_707_store_0_ack_0, ack => try1_CP_1680_elements(487)); -- 
    -- CP-element group 488:  transition  input  bypass 
    -- CP-element group 488: predecessors 
    -- CP-element group 488: 	390 
    -- CP-element group 488: successors 
    -- CP-element group 488: 	509 
    -- CP-element group 488:  members (5) 
      -- CP-element group 488: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_update_completed_
      -- CP-element group 488: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_Update/$exit
      -- CP-element group 488: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_Update/word_access_complete/$exit
      -- CP-element group 488: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_Update/word_access_complete/word_0/$exit
      -- CP-element group 488: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(488)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(488)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(488) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_707_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 488_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_707_store_0_ack_1, ack => try1_CP_1680_elements(488)); -- 
    -- CP-element group 489:  transition  input  bypass 
    -- CP-element group 489: predecessors 
    -- CP-element group 489: 	483 
    -- CP-element group 489: successors 
    -- CP-element group 489:  members (3) 
      -- CP-element group 489: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_714_sample_completed_
      -- CP-element group 489: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_714_Sample/$exit
      -- CP-element group 489: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_714_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(489)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(489)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(489) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_714_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 489_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_714_inst_ack_0, ack => try1_CP_1680_elements(489)); -- 
    -- CP-element group 490:  transition  input  bypass 
    -- CP-element group 490: predecessors 
    -- CP-element group 490: 	390 
    -- CP-element group 490: successors 
    -- CP-element group 490: 	491 
    -- CP-element group 490:  members (3) 
      -- CP-element group 490: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_714_update_completed_
      -- CP-element group 490: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_714_Update/$exit
      -- CP-element group 490: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_714_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(490)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(490)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(490) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_714_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 490_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_714_inst_ack_1, ack => try1_CP_1680_elements(490)); -- 
    -- CP-element group 491:  join  transition  output  bypass 
    -- CP-element group 491: predecessors 
    -- CP-element group 491: 	390 
    -- CP-element group 491: 	506 
    -- CP-element group 491: 	490 
    -- CP-element group 491: successors 
    -- CP-element group 491: 	492 
    -- CP-element group 491:  members (9) 
      -- CP-element group 491: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_sample_start_
      -- CP-element group 491: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_Sample/$entry
      -- CP-element group 491: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_Sample/array_obj_ref_712_Split/$entry
      -- CP-element group 491: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_Sample/array_obj_ref_712_Split/$exit
      -- CP-element group 491: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_Sample/array_obj_ref_712_Split/split_req
      -- CP-element group 491: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_Sample/array_obj_ref_712_Split/split_ack
      -- CP-element group 491: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_Sample/word_access_start/$entry
      -- CP-element group 491: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_Sample/word_access_start/word_0/$entry
      -- CP-element group 491: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(491)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(491)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(491) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_712_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(491), ack => array_obj_ref_712_store_0_req_0); -- 
    try1_cp_element_group_491: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_491"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(390) & try1_CP_1680_elements(506) & try1_CP_1680_elements(490);
      gj_try1_cp_element_group_491 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(491), clk => clk, reset => reset); --
    end block;
    -- CP-element group 492:  transition  input  bypass 
    -- CP-element group 492: predecessors 
    -- CP-element group 492: 	491 
    -- CP-element group 492: successors 
    -- CP-element group 492: 	507 
    -- CP-element group 492:  members (5) 
      -- CP-element group 492: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_sample_completed_
      -- CP-element group 492: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_Sample/$exit
      -- CP-element group 492: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_Sample/word_access_start/$exit
      -- CP-element group 492: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_Sample/word_access_start/word_0/$exit
      -- CP-element group 492: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(492)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(492)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(492) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_712_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 492_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_712_store_0_ack_0, ack => try1_CP_1680_elements(492)); -- 
    -- CP-element group 493:  transition  input  bypass 
    -- CP-element group 493: predecessors 
    -- CP-element group 493: 	390 
    -- CP-element group 493: successors 
    -- CP-element group 493: 	509 
    -- CP-element group 493:  members (5) 
      -- CP-element group 493: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_update_completed_
      -- CP-element group 493: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_Update/$exit
      -- CP-element group 493: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_Update/word_access_complete/$exit
      -- CP-element group 493: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_Update/word_access_complete/word_0/$exit
      -- CP-element group 493: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(493)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(493)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(493) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_712_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 493_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_712_store_0_ack_1, ack => try1_CP_1680_elements(493)); -- 
    -- CP-element group 494:  transition  input  bypass 
    -- CP-element group 494: predecessors 
    -- CP-element group 494: 	483 
    -- CP-element group 494: successors 
    -- CP-element group 494:  members (3) 
      -- CP-element group 494: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_719_sample_completed_
      -- CP-element group 494: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_719_Sample/$exit
      -- CP-element group 494: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_719_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(494)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(494)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(494) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_719_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 494_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_719_inst_ack_0, ack => try1_CP_1680_elements(494)); -- 
    -- CP-element group 495:  transition  input  bypass 
    -- CP-element group 495: predecessors 
    -- CP-element group 495: 	390 
    -- CP-element group 495: successors 
    -- CP-element group 495: 	496 
    -- CP-element group 495:  members (3) 
      -- CP-element group 495: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_719_update_completed_
      -- CP-element group 495: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_719_Update/$exit
      -- CP-element group 495: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_719_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(495)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(495)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(495) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_719_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 495_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_719_inst_ack_1, ack => try1_CP_1680_elements(495)); -- 
    -- CP-element group 496:  join  transition  output  bypass 
    -- CP-element group 496: predecessors 
    -- CP-element group 496: 	390 
    -- CP-element group 496: 	495 
    -- CP-element group 496: 	507 
    -- CP-element group 496: successors 
    -- CP-element group 496: 	497 
    -- CP-element group 496:  members (9) 
      -- CP-element group 496: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_sample_start_
      -- CP-element group 496: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_Sample/$entry
      -- CP-element group 496: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_Sample/array_obj_ref_717_Split/$entry
      -- CP-element group 496: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_Sample/array_obj_ref_717_Split/$exit
      -- CP-element group 496: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_Sample/array_obj_ref_717_Split/split_req
      -- CP-element group 496: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_Sample/array_obj_ref_717_Split/split_ack
      -- CP-element group 496: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_Sample/word_access_start/$entry
      -- CP-element group 496: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_Sample/word_access_start/word_0/$entry
      -- CP-element group 496: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(496)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(496)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(496) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_717_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(496), ack => array_obj_ref_717_store_0_req_0); -- 
    try1_cp_element_group_496: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_496"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(390) & try1_CP_1680_elements(495) & try1_CP_1680_elements(507);
      gj_try1_cp_element_group_496 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(496), clk => clk, reset => reset); --
    end block;
    -- CP-element group 497:  transition  input  bypass 
    -- CP-element group 497: predecessors 
    -- CP-element group 497: 	496 
    -- CP-element group 497: successors 
    -- CP-element group 497: 	508 
    -- CP-element group 497:  members (5) 
      -- CP-element group 497: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_sample_completed_
      -- CP-element group 497: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_Sample/$exit
      -- CP-element group 497: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_Sample/word_access_start/$exit
      -- CP-element group 497: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_Sample/word_access_start/word_0/$exit
      -- CP-element group 497: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(497)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(497)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(497) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_717_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 497_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_717_store_0_ack_0, ack => try1_CP_1680_elements(497)); -- 
    -- CP-element group 498:  transition  input  bypass 
    -- CP-element group 498: predecessors 
    -- CP-element group 498: 	390 
    -- CP-element group 498: successors 
    -- CP-element group 498: 	509 
    -- CP-element group 498:  members (5) 
      -- CP-element group 498: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_update_completed_
      -- CP-element group 498: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_Update/$exit
      -- CP-element group 498: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_Update/word_access_complete/$exit
      -- CP-element group 498: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_Update/word_access_complete/word_0/$exit
      -- CP-element group 498: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(498)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(498)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(498) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_717_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 498_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_717_store_0_ack_1, ack => try1_CP_1680_elements(498)); -- 
    -- CP-element group 499:  transition  input  bypass 
    -- CP-element group 499: predecessors 
    -- CP-element group 499: 	483 
    -- CP-element group 499: successors 
    -- CP-element group 499:  members (3) 
      -- CP-element group 499: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_724_sample_completed_
      -- CP-element group 499: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_724_Sample/$exit
      -- CP-element group 499: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_724_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(499)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(499)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(499) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_724_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 499_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_724_inst_ack_0, ack => try1_CP_1680_elements(499)); -- 
    -- CP-element group 500:  transition  input  bypass 
    -- CP-element group 500: predecessors 
    -- CP-element group 500: 	390 
    -- CP-element group 500: successors 
    -- CP-element group 500: 	501 
    -- CP-element group 500:  members (3) 
      -- CP-element group 500: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_724_update_completed_
      -- CP-element group 500: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_724_Update/$exit
      -- CP-element group 500: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/slice_724_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(500)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(500)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(500) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:slice_724_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 500_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_724_inst_ack_1, ack => try1_CP_1680_elements(500)); -- 
    -- CP-element group 501:  join  transition  output  bypass 
    -- CP-element group 501: predecessors 
    -- CP-element group 501: 	390 
    -- CP-element group 501: 	500 
    -- CP-element group 501: 	508 
    -- CP-element group 501: successors 
    -- CP-element group 501: 	502 
    -- CP-element group 501:  members (9) 
      -- CP-element group 501: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_sample_start_
      -- CP-element group 501: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_Sample/$entry
      -- CP-element group 501: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_Sample/array_obj_ref_722_Split/$entry
      -- CP-element group 501: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_Sample/array_obj_ref_722_Split/$exit
      -- CP-element group 501: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_Sample/array_obj_ref_722_Split/split_req
      -- CP-element group 501: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_Sample/array_obj_ref_722_Split/split_ack
      -- CP-element group 501: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_Sample/word_access_start/$entry
      -- CP-element group 501: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_Sample/word_access_start/word_0/$entry
      -- CP-element group 501: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group try1_CP_1680_elements(501)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(501)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(501) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_722_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(501), ack => array_obj_ref_722_store_0_req_0); -- 
    try1_cp_element_group_501: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_501"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try1_CP_1680_elements(390) & try1_CP_1680_elements(500) & try1_CP_1680_elements(508);
      gj_try1_cp_element_group_501 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(501), clk => clk, reset => reset); --
    end block;
    -- CP-element group 502:  transition  input  bypass 
    -- CP-element group 502: predecessors 
    -- CP-element group 502: 	501 
    -- CP-element group 502: successors 
    -- CP-element group 502:  members (5) 
      -- CP-element group 502: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_sample_completed_
      -- CP-element group 502: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_Sample/$exit
      -- CP-element group 502: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_Sample/word_access_start/$exit
      -- CP-element group 502: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_Sample/word_access_start/word_0/$exit
      -- CP-element group 502: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(502)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(502)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(502) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_722_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 502_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_722_store_0_ack_0, ack => try1_CP_1680_elements(502)); -- 
    -- CP-element group 503:  transition  input  bypass 
    -- CP-element group 503: predecessors 
    -- CP-element group 503: 	390 
    -- CP-element group 503: successors 
    -- CP-element group 503: 	509 
    -- CP-element group 503:  members (5) 
      -- CP-element group 503: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_update_completed_
      -- CP-element group 503: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_Update/$exit
      -- CP-element group 503: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_Update/word_access_complete/$exit
      -- CP-element group 503: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_Update/word_access_complete/word_0/$exit
      -- CP-element group 503: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_722_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(503)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(503)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(503) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:array_obj_ref_722_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 503_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_722_store_0_ack_1, ack => try1_CP_1680_elements(503)); -- 
    -- CP-element group 504:  transition  input  bypass 
    -- CP-element group 504: predecessors 
    -- CP-element group 504: 	390 
    -- CP-element group 504: successors 
    -- CP-element group 504:  members (3) 
      -- CP-element group 504: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_729_sample_completed_
      -- CP-element group 504: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_729_Sample/$exit
      -- CP-element group 504: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_729_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(504)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(504)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(504) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_729_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 504_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_729_inst_ack_0, ack => try1_CP_1680_elements(504)); -- 
    -- CP-element group 505:  transition  input  bypass 
    -- CP-element group 505: predecessors 
    -- CP-element group 505: 	390 
    -- CP-element group 505: successors 
    -- CP-element group 505: 	509 
    -- CP-element group 505:  members (3) 
      -- CP-element group 505: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_729_update_completed_
      -- CP-element group 505: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_729_Update/$exit
      -- CP-element group 505: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/ADD_u12_u12_729_Update/ca
      -- 
    -- logger for CP element group try1_CP_1680_elements(505)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(505)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(505) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_729_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 505_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_729_inst_ack_1, ack => try1_CP_1680_elements(505)); -- 
    -- CP-element group 506:  transition  delay-element  bypass 
    -- CP-element group 506: predecessors 
    -- CP-element group 506: 	487 
    -- CP-element group 506: successors 
    -- CP-element group 506: 	491 
    -- CP-element group 506:  members (1) 
      -- CP-element group 506: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_707_array_obj_ref_712_delay
      -- 
    -- logger for CP element group try1_CP_1680_elements(506)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(506)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(506) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(506) is a control-delay.
    cp_element_506_delay: control_delay_element  generic map(name => " 506_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(487), ack => try1_CP_1680_elements(506), clk => clk, reset =>reset);
    -- CP-element group 507:  transition  delay-element  bypass 
    -- CP-element group 507: predecessors 
    -- CP-element group 507: 	492 
    -- CP-element group 507: successors 
    -- CP-element group 507: 	496 
    -- CP-element group 507:  members (1) 
      -- CP-element group 507: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_712_array_obj_ref_717_delay
      -- 
    -- logger for CP element group try1_CP_1680_elements(507)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(507)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(507) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(507) is a control-delay.
    cp_element_507_delay: control_delay_element  generic map(name => " 507_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(492), ack => try1_CP_1680_elements(507), clk => clk, reset =>reset);
    -- CP-element group 508:  transition  delay-element  bypass 
    -- CP-element group 508: predecessors 
    -- CP-element group 508: 	497 
    -- CP-element group 508: successors 
    -- CP-element group 508: 	501 
    -- CP-element group 508:  members (1) 
      -- CP-element group 508: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/array_obj_ref_717_array_obj_ref_722_delay
      -- 
    -- logger for CP element group try1_CP_1680_elements(508)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(508)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(508) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group try1_CP_1680_elements(508) is a control-delay.
    cp_element_508_delay: control_delay_element  generic map(name => " 508_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(497), ack => try1_CP_1680_elements(508), clk => clk, reset =>reset);
    -- CP-element group 509:  branch  join  transition  place  output  bypass 
    -- CP-element group 509: predecessors 
    -- CP-element group 509: 	493 
    -- CP-element group 509: 	498 
    -- CP-element group 509: 	503 
    -- CP-element group 509: 	505 
    -- CP-element group 509: 	488 
    -- CP-element group 509: successors 
    -- CP-element group 509: 	510 
    -- CP-element group 509: 	511 
    -- CP-element group 509:  members (24) 
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730__exit__
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731__entry__
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/call_stmt_705_to_assign_stmt_730/$exit
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_dead_link/$entry
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_eval_test/$entry
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_eval_test/$exit
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_eval_test/ULT_u12_u1_734/$entry
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_eval_test/ULT_u12_u1_734/$exit
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_eval_test/ULT_u12_u1_734/ULT_u12_u1_734_inputs/$entry
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_eval_test/ULT_u12_u1_734/ULT_u12_u1_734_inputs/$exit
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_eval_test/ULT_u12_u1_734/SplitProtocol/$entry
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_eval_test/ULT_u12_u1_734/SplitProtocol/$exit
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_eval_test/ULT_u12_u1_734/SplitProtocol/Sample/$entry
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_eval_test/ULT_u12_u1_734/SplitProtocol/Sample/$exit
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_eval_test/ULT_u12_u1_734/SplitProtocol/Sample/rr
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_eval_test/ULT_u12_u1_734/SplitProtocol/Sample/ra
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_eval_test/ULT_u12_u1_734/SplitProtocol/Update/$entry
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_eval_test/ULT_u12_u1_734/SplitProtocol/Update/$exit
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_eval_test/ULT_u12_u1_734/SplitProtocol/Update/cr
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_eval_test/ULT_u12_u1_734/SplitProtocol/Update/ca
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_eval_test/branch_req
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/ULT_u12_u1_734_place
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_if_link/$entry
      -- CP-element group 509: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_else_link/$entry
      -- 
    -- logger for CP element group try1_CP_1680_elements(509)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(509)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(509) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:if_stmt_731_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    branch_req_4747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(509), ack => if_stmt_731_branch_req_0); -- 
    try1_cp_element_group_509: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_509"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= try1_CP_1680_elements(493) & try1_CP_1680_elements(498) & try1_CP_1680_elements(503) & try1_CP_1680_elements(505) & try1_CP_1680_elements(488);
      gj_try1_cp_element_group_509 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(509), clk => clk, reset => reset); --
    end block;
    -- CP-element group 510:  fork  transition  place  input  output  bypass 
    -- CP-element group 510: predecessors 
    -- CP-element group 510: 	509 
    -- CP-element group 510: successors 
    -- CP-element group 510: 	513 
    -- CP-element group 510: 	514 
    -- CP-element group 510:  members (11) 
      -- CP-element group 510: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_if_link/$exit
      -- CP-element group 510: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_if_link/if_choice_transition
      -- CP-element group 510: 	 branch_block_stmt_443/branch_block_stmt_565/loopback
      -- CP-element group 510: 	 branch_block_stmt_443/branch_block_stmt_565/loopback_PhiReq/$entry
      -- CP-element group 510: 	 branch_block_stmt_443/branch_block_stmt_565/loopback_PhiReq/phi_stmt_567/$entry
      -- CP-element group 510: 	 branch_block_stmt_443/branch_block_stmt_565/loopback_PhiReq/phi_stmt_567/phi_stmt_567_sources/$entry
      -- CP-element group 510: 	 branch_block_stmt_443/branch_block_stmt_565/loopback_PhiReq/phi_stmt_567/phi_stmt_567_sources/Interlock/$entry
      -- CP-element group 510: 	 branch_block_stmt_443/branch_block_stmt_565/loopback_PhiReq/phi_stmt_567/phi_stmt_567_sources/Interlock/Sample/$entry
      -- CP-element group 510: 	 branch_block_stmt_443/branch_block_stmt_565/loopback_PhiReq/phi_stmt_567/phi_stmt_567_sources/Interlock/Sample/req
      -- CP-element group 510: 	 branch_block_stmt_443/branch_block_stmt_565/loopback_PhiReq/phi_stmt_567/phi_stmt_567_sources/Interlock/Update/$entry
      -- CP-element group 510: 	 branch_block_stmt_443/branch_block_stmt_565/loopback_PhiReq/phi_stmt_567/phi_stmt_567_sources/Interlock/Update/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(510)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(510)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(510) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:if_stmt_731_branch_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NL_730_571_buf_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NL_730_571_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_4752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 510_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_731_branch_ack_1, ack => try1_CP_1680_elements(510)); -- 
    req_4788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(510), ack => NL_730_571_buf_req_0); -- 
    req_4793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(510), ack => NL_730_571_buf_req_1); -- 
    -- CP-element group 511:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 511: predecessors 
    -- CP-element group 511: 	509 
    -- CP-element group 511: successors 
    -- CP-element group 511: 	518 
    -- CP-element group 511: 	519 
    -- CP-element group 511:  members (14) 
      -- CP-element group 511: 	 branch_block_stmt_443/assign_stmt_742__entry__
      -- CP-element group 511: 	 branch_block_stmt_443/branch_block_stmt_565__exit__
      -- CP-element group 511: 	 branch_block_stmt_443/branch_block_stmt_565/branch_block_stmt_565__exit__
      -- CP-element group 511: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731__exit__
      -- CP-element group 511: 	 branch_block_stmt_443/branch_block_stmt_565/$exit
      -- CP-element group 511: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_else_link/$exit
      -- CP-element group 511: 	 branch_block_stmt_443/branch_block_stmt_565/if_stmt_731_else_link/else_choice_transition
      -- CP-element group 511: 	 branch_block_stmt_443/assign_stmt_742/$entry
      -- CP-element group 511: 	 branch_block_stmt_443/assign_stmt_742/ADD_u12_u12_741_sample_start_
      -- CP-element group 511: 	 branch_block_stmt_443/assign_stmt_742/ADD_u12_u12_741_update_start_
      -- CP-element group 511: 	 branch_block_stmt_443/assign_stmt_742/ADD_u12_u12_741_Sample/$entry
      -- CP-element group 511: 	 branch_block_stmt_443/assign_stmt_742/ADD_u12_u12_741_Sample/rr
      -- CP-element group 511: 	 branch_block_stmt_443/assign_stmt_742/ADD_u12_u12_741_Update/$entry
      -- CP-element group 511: 	 branch_block_stmt_443/assign_stmt_742/ADD_u12_u12_741_Update/cr
      -- 
    -- logger for CP element group try1_CP_1680_elements(511)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(511)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(511) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:if_stmt_731_branch_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_741_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_741_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_4756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 511_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_731_branch_ack_0, ack => try1_CP_1680_elements(511)); -- 
    rr_4811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(511), ack => ADD_u12_u12_741_inst_req_0); -- 
    cr_4816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(511), ack => ADD_u12_u12_741_inst_req_1); -- 
    -- CP-element group 512:  transition  output  delay-element  bypass 
    -- CP-element group 512: predecessors 
    -- CP-element group 512: 	131 
    -- CP-element group 512: successors 
    -- CP-element group 512: 	516 
    -- CP-element group 512:  members (5) 
      -- CP-element group 512: 	 branch_block_stmt_443/branch_block_stmt_565/merge_stmt_566__entry___PhiReq/$exit
      -- CP-element group 512: 	 branch_block_stmt_443/branch_block_stmt_565/merge_stmt_566__entry___PhiReq/phi_stmt_567/$exit
      -- CP-element group 512: 	 branch_block_stmt_443/branch_block_stmt_565/merge_stmt_566__entry___PhiReq/phi_stmt_567/phi_stmt_567_sources/$exit
      -- CP-element group 512: 	 branch_block_stmt_443/branch_block_stmt_565/merge_stmt_566__entry___PhiReq/phi_stmt_567/phi_stmt_567_sources/type_cast_570_konst_delay_trans
      -- CP-element group 512: 	 branch_block_stmt_443/branch_block_stmt_565/merge_stmt_566__entry___PhiReq/phi_stmt_567/phi_stmt_567_req
      -- 
    -- logger for CP element group try1_CP_1680_elements(512)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(512)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(512) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:phi_stmt_567_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_567_req_4772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_567_req_4772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(512), ack => phi_stmt_567_req_0); -- 
    -- Element group try1_CP_1680_elements(512) is a control-delay.
    cp_element_512_delay: control_delay_element  generic map(name => " 512_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(131), ack => try1_CP_1680_elements(512), clk => clk, reset =>reset);
    -- CP-element group 513:  transition  input  bypass 
    -- CP-element group 513: predecessors 
    -- CP-element group 513: 	510 
    -- CP-element group 513: successors 
    -- CP-element group 513: 	515 
    -- CP-element group 513:  members (2) 
      -- CP-element group 513: 	 branch_block_stmt_443/branch_block_stmt_565/loopback_PhiReq/phi_stmt_567/phi_stmt_567_sources/Interlock/Sample/$exit
      -- CP-element group 513: 	 branch_block_stmt_443/branch_block_stmt_565/loopback_PhiReq/phi_stmt_567/phi_stmt_567_sources/Interlock/Sample/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(513)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(513)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(513) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NL_730_571_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 513_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NL_730_571_buf_ack_0, ack => try1_CP_1680_elements(513)); -- 
    -- CP-element group 514:  transition  input  bypass 
    -- CP-element group 514: predecessors 
    -- CP-element group 514: 	510 
    -- CP-element group 514: successors 
    -- CP-element group 514: 	515 
    -- CP-element group 514:  members (2) 
      -- CP-element group 514: 	 branch_block_stmt_443/branch_block_stmt_565/loopback_PhiReq/phi_stmt_567/phi_stmt_567_sources/Interlock/Update/$exit
      -- CP-element group 514: 	 branch_block_stmt_443/branch_block_stmt_565/loopback_PhiReq/phi_stmt_567/phi_stmt_567_sources/Interlock/Update/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(514)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(514)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(514) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NL_730_571_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_4794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 514_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NL_730_571_buf_ack_1, ack => try1_CP_1680_elements(514)); -- 
    -- CP-element group 515:  join  transition  output  bypass 
    -- CP-element group 515: predecessors 
    -- CP-element group 515: 	513 
    -- CP-element group 515: 	514 
    -- CP-element group 515: successors 
    -- CP-element group 515: 	516 
    -- CP-element group 515:  members (5) 
      -- CP-element group 515: 	 branch_block_stmt_443/branch_block_stmt_565/loopback_PhiReq/$exit
      -- CP-element group 515: 	 branch_block_stmt_443/branch_block_stmt_565/loopback_PhiReq/phi_stmt_567/$exit
      -- CP-element group 515: 	 branch_block_stmt_443/branch_block_stmt_565/loopback_PhiReq/phi_stmt_567/phi_stmt_567_sources/$exit
      -- CP-element group 515: 	 branch_block_stmt_443/branch_block_stmt_565/loopback_PhiReq/phi_stmt_567/phi_stmt_567_sources/Interlock/$exit
      -- CP-element group 515: 	 branch_block_stmt_443/branch_block_stmt_565/loopback_PhiReq/phi_stmt_567/phi_stmt_567_req
      -- 
    -- logger for CP element group try1_CP_1680_elements(515)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(515)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(515) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:phi_stmt_567_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_567_req_4795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_567_req_4795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(515), ack => phi_stmt_567_req_1); -- 
    try1_cp_element_group_515: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_515"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(513) & try1_CP_1680_elements(514);
      gj_try1_cp_element_group_515 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(515), clk => clk, reset => reset); --
    end block;
    -- CP-element group 516:  merge  transition  place  bypass 
    -- CP-element group 516: predecessors 
    -- CP-element group 516: 	512 
    -- CP-element group 516: 	515 
    -- CP-element group 516: successors 
    -- CP-element group 516: 	517 
    -- CP-element group 516:  members (2) 
      -- CP-element group 516: 	 branch_block_stmt_443/branch_block_stmt_565/merge_stmt_566_PhiReqMerge
      -- CP-element group 516: 	 branch_block_stmt_443/branch_block_stmt_565/merge_stmt_566_PhiAck/$entry
      -- 
    -- logger for CP element group try1_CP_1680_elements(516)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(516)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(516) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(516) <= OrReduce(try1_CP_1680_elements(512) & try1_CP_1680_elements(515));
    -- CP-element group 517:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 517: predecessors 
    -- CP-element group 517: 	516 
    -- CP-element group 517: successors 
    -- CP-element group 517: 	292 
    -- CP-element group 517: 	293 
    -- CP-element group 517:  members (21) 
      -- CP-element group 517: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575__entry__
      -- CP-element group 517: 	 branch_block_stmt_443/branch_block_stmt_565/merge_stmt_566__exit__
      -- CP-element group 517: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/$entry
      -- CP-element group 517: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_sample_start_
      -- CP-element group 517: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_update_start_
      -- CP-element group 517: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_word_address_calculated
      -- CP-element group 517: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_root_address_calculated
      -- CP-element group 517: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_Sample/$entry
      -- CP-element group 517: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_Sample/STORE_total_573_Split/$entry
      -- CP-element group 517: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_Sample/STORE_total_573_Split/$exit
      -- CP-element group 517: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_Sample/STORE_total_573_Split/split_req
      -- CP-element group 517: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_Sample/STORE_total_573_Split/split_ack
      -- CP-element group 517: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_Sample/word_access_start/$entry
      -- CP-element group 517: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_Sample/word_access_start/word_0/$entry
      -- CP-element group 517: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_Sample/word_access_start/word_0/rr
      -- CP-element group 517: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_Update/$entry
      -- CP-element group 517: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_Update/word_access_complete/$entry
      -- CP-element group 517: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_Update/word_access_complete/word_0/$entry
      -- CP-element group 517: 	 branch_block_stmt_443/branch_block_stmt_565/assign_stmt_575/STORE_total_573_Update/word_access_complete/word_0/cr
      -- CP-element group 517: 	 branch_block_stmt_443/branch_block_stmt_565/merge_stmt_566_PhiAck/$exit
      -- CP-element group 517: 	 branch_block_stmt_443/branch_block_stmt_565/merge_stmt_566_PhiAck/phi_stmt_567_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(517)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(517)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(517) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:phi_stmt_567_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:STORE_total_573_store_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:STORE_total_573_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_567_ack_4800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 517_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_567_ack_0, ack => try1_CP_1680_elements(517)); -- 
    rr_3251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(517), ack => STORE_total_573_store_0_req_0); -- 
    cr_3262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(517), ack => STORE_total_573_store_0_req_1); -- 
    -- CP-element group 518:  transition  input  bypass 
    -- CP-element group 518: predecessors 
    -- CP-element group 518: 	511 
    -- CP-element group 518: successors 
    -- CP-element group 518:  members (3) 
      -- CP-element group 518: 	 branch_block_stmt_443/assign_stmt_742/ADD_u12_u12_741_sample_completed_
      -- CP-element group 518: 	 branch_block_stmt_443/assign_stmt_742/ADD_u12_u12_741_Sample/$exit
      -- CP-element group 518: 	 branch_block_stmt_443/assign_stmt_742/ADD_u12_u12_741_Sample/ra
      -- 
    -- logger for CP element group try1_CP_1680_elements(518)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(518)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(518) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_741_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 518_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_741_inst_ack_0, ack => try1_CP_1680_elements(518)); -- 
    -- CP-element group 519:  branch  transition  place  input  output  bypass 
    -- CP-element group 519: predecessors 
    -- CP-element group 519: 	511 
    -- CP-element group 519: successors 
    -- CP-element group 519: 	520 
    -- CP-element group 519: 	521 
    -- CP-element group 519:  members (27) 
      -- CP-element group 519: 	 branch_block_stmt_443/assign_stmt_742__exit__
      -- CP-element group 519: 	 branch_block_stmt_443/if_stmt_743__entry__
      -- CP-element group 519: 	 branch_block_stmt_443/assign_stmt_742/$exit
      -- CP-element group 519: 	 branch_block_stmt_443/assign_stmt_742/ADD_u12_u12_741_update_completed_
      -- CP-element group 519: 	 branch_block_stmt_443/assign_stmt_742/ADD_u12_u12_741_Update/$exit
      -- CP-element group 519: 	 branch_block_stmt_443/assign_stmt_742/ADD_u12_u12_741_Update/ca
      -- CP-element group 519: 	 branch_block_stmt_443/if_stmt_743_dead_link/$entry
      -- CP-element group 519: 	 branch_block_stmt_443/if_stmt_743_eval_test/$entry
      -- CP-element group 519: 	 branch_block_stmt_443/if_stmt_743_eval_test/$exit
      -- CP-element group 519: 	 branch_block_stmt_443/if_stmt_743_eval_test/ULT_u12_u1_746/$entry
      -- CP-element group 519: 	 branch_block_stmt_443/if_stmt_743_eval_test/ULT_u12_u1_746/$exit
      -- CP-element group 519: 	 branch_block_stmt_443/if_stmt_743_eval_test/ULT_u12_u1_746/ULT_u12_u1_746_inputs/$entry
      -- CP-element group 519: 	 branch_block_stmt_443/if_stmt_743_eval_test/ULT_u12_u1_746/ULT_u12_u1_746_inputs/$exit
      -- CP-element group 519: 	 branch_block_stmt_443/if_stmt_743_eval_test/ULT_u12_u1_746/SplitProtocol/$entry
      -- CP-element group 519: 	 branch_block_stmt_443/if_stmt_743_eval_test/ULT_u12_u1_746/SplitProtocol/$exit
      -- CP-element group 519: 	 branch_block_stmt_443/if_stmt_743_eval_test/ULT_u12_u1_746/SplitProtocol/Sample/$entry
      -- CP-element group 519: 	 branch_block_stmt_443/if_stmt_743_eval_test/ULT_u12_u1_746/SplitProtocol/Sample/$exit
      -- CP-element group 519: 	 branch_block_stmt_443/if_stmt_743_eval_test/ULT_u12_u1_746/SplitProtocol/Sample/rr
      -- CP-element group 519: 	 branch_block_stmt_443/if_stmt_743_eval_test/ULT_u12_u1_746/SplitProtocol/Sample/ra
      -- CP-element group 519: 	 branch_block_stmt_443/if_stmt_743_eval_test/ULT_u12_u1_746/SplitProtocol/Update/$entry
      -- CP-element group 519: 	 branch_block_stmt_443/if_stmt_743_eval_test/ULT_u12_u1_746/SplitProtocol/Update/$exit
      -- CP-element group 519: 	 branch_block_stmt_443/if_stmt_743_eval_test/ULT_u12_u1_746/SplitProtocol/Update/cr
      -- CP-element group 519: 	 branch_block_stmt_443/if_stmt_743_eval_test/ULT_u12_u1_746/SplitProtocol/Update/ca
      -- CP-element group 519: 	 branch_block_stmt_443/if_stmt_743_eval_test/branch_req
      -- CP-element group 519: 	 branch_block_stmt_443/ULT_u12_u1_746_place
      -- CP-element group 519: 	 branch_block_stmt_443/if_stmt_743_if_link/$entry
      -- CP-element group 519: 	 branch_block_stmt_443/if_stmt_743_else_link/$entry
      -- 
    -- logger for CP element group try1_CP_1680_elements(519)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(519)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(519) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:ADD_u12_u12_741_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:if_stmt_743_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_4817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 519_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u12_u12_741_inst_ack_1, ack => try1_CP_1680_elements(519)); -- 
    branch_req_4844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(519), ack => if_stmt_743_branch_req_0); -- 
    -- CP-element group 520:  fork  transition  place  input  output  bypass 
    -- CP-element group 520: predecessors 
    -- CP-element group 520: 	519 
    -- CP-element group 520: successors 
    -- CP-element group 520: 	523 
    -- CP-element group 520: 	524 
    -- CP-element group 520:  members (11) 
      -- CP-element group 520: 	 branch_block_stmt_443/if_stmt_743_if_link/$exit
      -- CP-element group 520: 	 branch_block_stmt_443/if_stmt_743_if_link/if_choice_transition
      -- CP-element group 520: 	 branch_block_stmt_443/loopback
      -- CP-element group 520: 	 branch_block_stmt_443/loopback_PhiReq/$entry
      -- CP-element group 520: 	 branch_block_stmt_443/loopback_PhiReq/phi_stmt_445/$entry
      -- CP-element group 520: 	 branch_block_stmt_443/loopback_PhiReq/phi_stmt_445/phi_stmt_445_sources/$entry
      -- CP-element group 520: 	 branch_block_stmt_443/loopback_PhiReq/phi_stmt_445/phi_stmt_445_sources/Interlock/$entry
      -- CP-element group 520: 	 branch_block_stmt_443/loopback_PhiReq/phi_stmt_445/phi_stmt_445_sources/Interlock/Sample/$entry
      -- CP-element group 520: 	 branch_block_stmt_443/loopback_PhiReq/phi_stmt_445/phi_stmt_445_sources/Interlock/Sample/req
      -- CP-element group 520: 	 branch_block_stmt_443/loopback_PhiReq/phi_stmt_445/phi_stmt_445_sources/Interlock/Update/$entry
      -- CP-element group 520: 	 branch_block_stmt_443/loopback_PhiReq/phi_stmt_445/phi_stmt_445_sources/Interlock/Update/req
      -- 
    -- logger for CP element group try1_CP_1680_elements(520)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(520)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(520) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:if_stmt_743_branch_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NG_742_449_buf_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NG_742_449_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_4849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 520_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_743_branch_ack_1, ack => try1_CP_1680_elements(520)); -- 
    req_4885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(520), ack => NG_742_449_buf_req_0); -- 
    req_4890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(520), ack => NG_742_449_buf_req_1); -- 
    -- CP-element group 521:  merge  transition  place  input  bypass 
    -- CP-element group 521: predecessors 
    -- CP-element group 521: 	519 
    -- CP-element group 521: successors 
    -- CP-element group 521:  members (6) 
      -- CP-element group 521: 	 branch_block_stmt_443/branch_block_stmt_443__exit__
      -- CP-element group 521: 	 $exit
      -- CP-element group 521: 	 branch_block_stmt_443/if_stmt_743__exit__
      -- CP-element group 521: 	 branch_block_stmt_443/$exit
      -- CP-element group 521: 	 branch_block_stmt_443/if_stmt_743_else_link/$exit
      -- CP-element group 521: 	 branch_block_stmt_443/if_stmt_743_else_link/else_choice_transition
      -- 
    -- logger for CP element group try1_CP_1680_elements(521)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(521)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(521) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:if_stmt_743_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_4853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 521_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_743_branch_ack_0, ack => try1_CP_1680_elements(521)); -- 
    -- CP-element group 522:  transition  output  delay-element  bypass 
    -- CP-element group 522: predecessors 
    -- CP-element group 522: 	1 
    -- CP-element group 522: successors 
    -- CP-element group 522: 	526 
    -- CP-element group 522:  members (5) 
      -- CP-element group 522: 	 branch_block_stmt_443/merge_stmt_444__entry___PhiReq/$exit
      -- CP-element group 522: 	 branch_block_stmt_443/merge_stmt_444__entry___PhiReq/phi_stmt_445/$exit
      -- CP-element group 522: 	 branch_block_stmt_443/merge_stmt_444__entry___PhiReq/phi_stmt_445/phi_stmt_445_sources/$exit
      -- CP-element group 522: 	 branch_block_stmt_443/merge_stmt_444__entry___PhiReq/phi_stmt_445/phi_stmt_445_sources/type_cast_448_konst_delay_trans
      -- CP-element group 522: 	 branch_block_stmt_443/merge_stmt_444__entry___PhiReq/phi_stmt_445/phi_stmt_445_req
      -- 
    -- logger for CP element group try1_CP_1680_elements(522)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(522)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(522) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:phi_stmt_445_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_445_req_4869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_445_req_4869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(522), ack => phi_stmt_445_req_0); -- 
    -- Element group try1_CP_1680_elements(522) is a control-delay.
    cp_element_522_delay: control_delay_element  generic map(name => " 522_delay", delay_value => 1)  port map(req => try1_CP_1680_elements(1), ack => try1_CP_1680_elements(522), clk => clk, reset =>reset);
    -- CP-element group 523:  transition  input  bypass 
    -- CP-element group 523: predecessors 
    -- CP-element group 523: 	520 
    -- CP-element group 523: successors 
    -- CP-element group 523: 	525 
    -- CP-element group 523:  members (2) 
      -- CP-element group 523: 	 branch_block_stmt_443/loopback_PhiReq/phi_stmt_445/phi_stmt_445_sources/Interlock/Sample/$exit
      -- CP-element group 523: 	 branch_block_stmt_443/loopback_PhiReq/phi_stmt_445/phi_stmt_445_sources/Interlock/Sample/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(523)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(523)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(523) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NG_742_449_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 523_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NG_742_449_buf_ack_0, ack => try1_CP_1680_elements(523)); -- 
    -- CP-element group 524:  transition  input  bypass 
    -- CP-element group 524: predecessors 
    -- CP-element group 524: 	520 
    -- CP-element group 524: successors 
    -- CP-element group 524: 	525 
    -- CP-element group 524:  members (2) 
      -- CP-element group 524: 	 branch_block_stmt_443/loopback_PhiReq/phi_stmt_445/phi_stmt_445_sources/Interlock/Update/$exit
      -- CP-element group 524: 	 branch_block_stmt_443/loopback_PhiReq/phi_stmt_445/phi_stmt_445_sources/Interlock/Update/ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(524)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(524)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(524) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:NG_742_449_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_4891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 524_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NG_742_449_buf_ack_1, ack => try1_CP_1680_elements(524)); -- 
    -- CP-element group 525:  join  transition  output  bypass 
    -- CP-element group 525: predecessors 
    -- CP-element group 525: 	523 
    -- CP-element group 525: 	524 
    -- CP-element group 525: successors 
    -- CP-element group 525: 	526 
    -- CP-element group 525:  members (5) 
      -- CP-element group 525: 	 branch_block_stmt_443/loopback_PhiReq/$exit
      -- CP-element group 525: 	 branch_block_stmt_443/loopback_PhiReq/phi_stmt_445/$exit
      -- CP-element group 525: 	 branch_block_stmt_443/loopback_PhiReq/phi_stmt_445/phi_stmt_445_sources/$exit
      -- CP-element group 525: 	 branch_block_stmt_443/loopback_PhiReq/phi_stmt_445/phi_stmt_445_sources/Interlock/$exit
      -- CP-element group 525: 	 branch_block_stmt_443/loopback_PhiReq/phi_stmt_445/phi_stmt_445_req
      -- 
    -- logger for CP element group try1_CP_1680_elements(525)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(525)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(525) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:phi_stmt_445_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_445_req_4892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_445_req_4892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(525), ack => phi_stmt_445_req_1); -- 
    try1_cp_element_group_525: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "try1_cp_element_group_525"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_1680_elements(523) & try1_CP_1680_elements(524);
      gj_try1_cp_element_group_525 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_1680_elements(525), clk => clk, reset => reset); --
    end block;
    -- CP-element group 526:  merge  transition  place  bypass 
    -- CP-element group 526: predecessors 
    -- CP-element group 526: 	522 
    -- CP-element group 526: 	525 
    -- CP-element group 526: successors 
    -- CP-element group 526: 	527 
    -- CP-element group 526:  members (2) 
      -- CP-element group 526: 	 branch_block_stmt_443/merge_stmt_444_PhiReqMerge
      -- CP-element group 526: 	 branch_block_stmt_443/merge_stmt_444_PhiAck/$entry
      -- 
    -- logger for CP element group try1_CP_1680_elements(526)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(526)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(526) fired."); 
        -- 
      end if; --
    end process; 
    try1_CP_1680_elements(526) <= OrReduce(try1_CP_1680_elements(522) & try1_CP_1680_elements(525));
    -- CP-element group 527:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 527: predecessors 
    -- CP-element group 527: 	526 
    -- CP-element group 527: successors 
    -- CP-element group 527: 	129 
    -- CP-element group 527: 	130 
    -- CP-element group 527:  members (21) 
      -- CP-element group 527: 	 branch_block_stmt_443/merge_stmt_444__exit__
      -- CP-element group 527: 	 branch_block_stmt_443/assign_stmt_453__entry__
      -- CP-element group 527: 	 branch_block_stmt_443/assign_stmt_453/$entry
      -- CP-element group 527: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_sample_start_
      -- CP-element group 527: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_update_start_
      -- CP-element group 527: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_word_address_calculated
      -- CP-element group 527: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_root_address_calculated
      -- CP-element group 527: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_Sample/$entry
      -- CP-element group 527: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_Sample/STORE_PJ_451_Split/$entry
      -- CP-element group 527: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_Sample/STORE_PJ_451_Split/$exit
      -- CP-element group 527: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_Sample/STORE_PJ_451_Split/split_req
      -- CP-element group 527: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_Sample/STORE_PJ_451_Split/split_ack
      -- CP-element group 527: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_Sample/word_access_start/$entry
      -- CP-element group 527: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_Sample/word_access_start/word_0/$entry
      -- CP-element group 527: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_Sample/word_access_start/word_0/rr
      -- CP-element group 527: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_Update/$entry
      -- CP-element group 527: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_Update/word_access_complete/$entry
      -- CP-element group 527: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_Update/word_access_complete/word_0/$entry
      -- CP-element group 527: 	 branch_block_stmt_443/assign_stmt_453/STORE_PJ_451_Update/word_access_complete/word_0/cr
      -- CP-element group 527: 	 branch_block_stmt_443/merge_stmt_444_PhiAck/$exit
      -- CP-element group 527: 	 branch_block_stmt_443/merge_stmt_444_PhiAck/phi_stmt_445_ack
      -- 
    -- logger for CP element group try1_CP_1680_elements(527)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and try1_CP_1680_elements(527)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:try1_CP_1680_elements(527) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:phi_stmt_445_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:STORE_PJ_451_store_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:try1:CP:STORE_PJ_451_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_445_ack_4897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 527_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_445_ack_0, ack => try1_CP_1680_elements(527)); -- 
    rr_2360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(527), ack => STORE_PJ_451_store_0_req_0); -- 
    cr_2371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_1680_elements(527), ack => STORE_PJ_451_store_0_req_1); -- 
    try1_do_while_stmt_344_terminator_2319: loop_terminator -- 
      generic map (name => " try1_do_while_stmt_344_terminator_2319", max_iterations_in_flight =>7) 
      port map(loop_body_exit => try1_CP_1680_elements(6),loop_continue => try1_CP_1680_elements(127),loop_terminate => try1_CP_1680_elements(126),loop_back => try1_CP_1680_elements(4),loop_exit => try1_CP_1680_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_346_phi_seq_1753_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= try1_CP_1680_elements(18);
      try1_CP_1680_elements(21)<= src_sample_reqs(0);
      src_sample_acks(0)  <= try1_CP_1680_elements(21);
      try1_CP_1680_elements(22)<= src_update_reqs(0);
      src_update_acks(0)  <= try1_CP_1680_elements(23);
      try1_CP_1680_elements(19) <= phi_mux_reqs(0);
      triggers(1)  <= try1_CP_1680_elements(16);
      try1_CP_1680_elements(25)<= src_sample_reqs(1);
      src_sample_acks(1)  <= try1_CP_1680_elements(27);
      try1_CP_1680_elements(26)<= src_update_reqs(1);
      src_update_acks(1)  <= try1_CP_1680_elements(28);
      try1_CP_1680_elements(17) <= phi_mux_reqs(1);
      phi_stmt_346_phi_seq_1753 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_346_phi_seq_1753") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => try1_CP_1680_elements(11), 
          phi_sample_ack => try1_CP_1680_elements(14), 
          phi_update_req => try1_CP_1680_elements(13), 
          phi_update_ack => try1_CP_1680_elements(15), 
          phi_mux_ack => try1_CP_1680_elements(20), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1705_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= try1_CP_1680_elements(7);
        preds(1)  <= try1_CP_1680_elements(8);
        entry_tmerge_1705 : transition_merge -- 
          generic map(name => " entry_tmerge_1705")
          port map (preds => preds, symbol_out => try1_CP_1680_elements(9));
          -- 
    end block;
    try1_do_while_stmt_455_terminator_3208: loop_terminator -- 
      generic map (name => " try1_do_while_stmt_455_terminator_3208", max_iterations_in_flight =>7) 
      port map(loop_body_exit => try1_CP_1680_elements(136),loop_continue => try1_CP_1680_elements(290),loop_terminate => try1_CP_1680_elements(289),loop_back => try1_CP_1680_elements(134),loop_exit => try1_CP_1680_elements(133),clk => clk, reset => reset); -- 
    phi_stmt_457_phi_seq_2443_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= try1_CP_1680_elements(148);
      try1_CP_1680_elements(151)<= src_sample_reqs(0);
      src_sample_acks(0)  <= try1_CP_1680_elements(151);
      try1_CP_1680_elements(152)<= src_update_reqs(0);
      src_update_acks(0)  <= try1_CP_1680_elements(153);
      try1_CP_1680_elements(149) <= phi_mux_reqs(0);
      triggers(1)  <= try1_CP_1680_elements(146);
      try1_CP_1680_elements(155)<= src_sample_reqs(1);
      src_sample_acks(1)  <= try1_CP_1680_elements(157);
      try1_CP_1680_elements(156)<= src_update_reqs(1);
      src_update_acks(1)  <= try1_CP_1680_elements(158);
      try1_CP_1680_elements(147) <= phi_mux_reqs(1);
      phi_stmt_457_phi_seq_2443 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_457_phi_seq_2443") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => try1_CP_1680_elements(141), 
          phi_sample_ack => try1_CP_1680_elements(144), 
          phi_update_req => try1_CP_1680_elements(143), 
          phi_update_ack => try1_CP_1680_elements(145), 
          phi_mux_ack => try1_CP_1680_elements(150), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2395_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= try1_CP_1680_elements(137);
        preds(1)  <= try1_CP_1680_elements(138);
        entry_tmerge_2395 : transition_merge -- 
          generic map(name => " entry_tmerge_2395")
          port map (preds => preds, symbol_out => try1_CP_1680_elements(139));
          -- 
    end block;
    try1_do_while_stmt_577_terminator_3721: loop_terminator -- 
      generic map (name => " try1_do_while_stmt_577_terminator_3721", max_iterations_in_flight =>7) 
      port map(loop_body_exit => try1_CP_1680_elements(299),loop_continue => try1_CP_1680_elements(368),loop_terminate => try1_CP_1680_elements(367),loop_back => try1_CP_1680_elements(297),loop_exit => try1_CP_1680_elements(296),clk => clk, reset => reset); -- 
    phi_stmt_579_phi_seq_3334_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= try1_CP_1680_elements(311);
      try1_CP_1680_elements(314)<= src_sample_reqs(0);
      src_sample_acks(0)  <= try1_CP_1680_elements(314);
      try1_CP_1680_elements(315)<= src_update_reqs(0);
      src_update_acks(0)  <= try1_CP_1680_elements(316);
      try1_CP_1680_elements(312) <= phi_mux_reqs(0);
      triggers(1)  <= try1_CP_1680_elements(309);
      try1_CP_1680_elements(318)<= src_sample_reqs(1);
      src_sample_acks(1)  <= try1_CP_1680_elements(320);
      try1_CP_1680_elements(319)<= src_update_reqs(1);
      src_update_acks(1)  <= try1_CP_1680_elements(321);
      try1_CP_1680_elements(310) <= phi_mux_reqs(1);
      phi_stmt_579_phi_seq_3334 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_579_phi_seq_3334") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => try1_CP_1680_elements(304), 
          phi_sample_ack => try1_CP_1680_elements(307), 
          phi_update_req => try1_CP_1680_elements(306), 
          phi_update_ack => try1_CP_1680_elements(308), 
          phi_mux_ack => try1_CP_1680_elements(313), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3286_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= try1_CP_1680_elements(300);
        preds(1)  <= try1_CP_1680_elements(301);
        entry_tmerge_3286 : transition_merge -- 
          generic map(name => " entry_tmerge_3286")
          port map (preds => preds, symbol_out => try1_CP_1680_elements(302));
          -- 
    end block;
    try1_do_while_stmt_640_terminator_4484: loop_terminator -- 
      generic map (name => " try1_do_while_stmt_640_terminator_4484", max_iterations_in_flight =>7) 
      port map(loop_body_exit => try1_CP_1680_elements(395),loop_continue => try1_CP_1680_elements(478),loop_terminate => try1_CP_1680_elements(477),loop_back => try1_CP_1680_elements(393),loop_exit => try1_CP_1680_elements(392),clk => clk, reset => reset); -- 
    phi_stmt_642_phi_seq_3995_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= try1_CP_1680_elements(407);
      try1_CP_1680_elements(410)<= src_sample_reqs(0);
      src_sample_acks(0)  <= try1_CP_1680_elements(410);
      try1_CP_1680_elements(411)<= src_update_reqs(0);
      src_update_acks(0)  <= try1_CP_1680_elements(412);
      try1_CP_1680_elements(408) <= phi_mux_reqs(0);
      triggers(1)  <= try1_CP_1680_elements(405);
      try1_CP_1680_elements(414)<= src_sample_reqs(1);
      src_sample_acks(1)  <= try1_CP_1680_elements(416);
      try1_CP_1680_elements(415)<= src_update_reqs(1);
      src_update_acks(1)  <= try1_CP_1680_elements(417);
      try1_CP_1680_elements(406) <= phi_mux_reqs(1);
      phi_stmt_642_phi_seq_3995 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_642_phi_seq_3995") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => try1_CP_1680_elements(400), 
          phi_sample_ack => try1_CP_1680_elements(403), 
          phi_update_req => try1_CP_1680_elements(402), 
          phi_update_ack => try1_CP_1680_elements(404), 
          phi_mux_ack => try1_CP_1680_elements(409), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3947_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= try1_CP_1680_elements(396);
        preds(1)  <= try1_CP_1680_elements(397);
        entry_tmerge_3947 : transition_merge -- 
          generic map(name => " entry_tmerge_3947")
          port map (preds => preds, symbol_out => try1_CP_1680_elements(398));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u12_u12_621_wire : std_logic_vector(11 downto 0);
    signal ADD_u12_u12_629_wire : std_logic_vector(11 downto 0);
    signal ADD_u12_u12_700_wire : std_logic_vector(11 downto 0);
    signal ADD_u12_u12_702_wire : std_logic_vector(11 downto 0);
    signal ADD_u16_u16_558_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_606_wire : std_logic_vector(15 downto 0);
    signal G_445 : std_logic_vector(11 downto 0);
    signal HHHH_678 : std_logic_vector(11 downto 0);
    signal HHH_594_delayed_4_0_681 : std_logic_vector(11 downto 0);
    signal HHH_665 : std_logic_vector(11 downto 0);
    signal HH_584_delayed_4_0_668 : std_logic_vector(11 downto 0);
    signal HH_652 : std_logic_vector(11 downto 0);
    signal H_574_delayed_5_0_655 : std_logic_vector(11 downto 0);
    signal H_642 : std_logic_vector(11 downto 0);
    signal J_457 : std_logic_vector(11 downto 0);
    signal K_517_delayed_5_0_595 : std_logic_vector(31 downto 0);
    signal K_579 : std_logic_vector(31 downto 0);
    signal LOAD_PJ_500_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_PJ_500_wire : std_logic_vector(15 downto 0);
    signal LOAD_PJ_500_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_PJ_505_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_PJ_505_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_PJ_527_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_PJ_527_wire : std_logic_vector(15 downto 0);
    signal LOAD_PJ_527_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_PJ_532_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_PJ_532_wire : std_logic_vector(15 downto 0);
    signal LOAD_PJ_532_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_PJ_556_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_PJ_556_wire : std_logic_vector(15 downto 0);
    signal LOAD_PJ_556_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_ZJ_357_data_0 : std_logic_vector(11 downto 0);
    signal LOAD_ZJ_357_wire : std_logic_vector(11 downto 0);
    signal LOAD_ZJ_357_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_one_366_data_0 : std_logic_vector(0 downto 0);
    signal LOAD_one_366_wire : std_logic_vector(0 downto 0);
    signal LOAD_one_366_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_one_475_data_0 : std_logic_vector(0 downto 0);
    signal LOAD_one_475_wire : std_logic_vector(0 downto 0);
    signal LOAD_one_475_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_total_603_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_total_603_wire : std_logic_vector(15 downto 0);
    signal LOAD_total_603_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_total_622_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_total_622_wire : std_logic_vector(15 downto 0);
    signal LOAD_total_622_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_zer_626_data_0 : std_logic_vector(3 downto 0);
    signal LOAD_zer_626_wire : std_logic_vector(3 downto 0);
    signal LOAD_zer_626_word_address_0 : std_logic_vector(0 downto 0);
    signal L_567 : std_logic_vector(11 downto 0);
    signal MUL_u16_u16_600_wire : std_logic_vector(15 downto 0);
    signal NGG_420_delayed_4_0_481 : std_logic_vector(31 downto 0);
    signal NGG_470 : std_logic_vector(31 downto 0);
    signal NG_742 : std_logic_vector(11 downto 0);
    signal NG_742_449_buffered : std_logic_vector(11 downto 0);
    signal NH_691 : std_logic_vector(11 downto 0);
    signal NH_691_646_buffered : std_logic_vector(11 downto 0);
    signal NJJ_415_delayed_2_0_473 : std_logic_vector(30 downto 0);
    signal NJJ_466 : std_logic_vector(30 downto 0);
    signal NJ_554 : std_logic_vector(11 downto 0);
    signal NJ_554_461_buffered : std_logic_vector(11 downto 0);
    signal NK_612 : std_logic_vector(31 downto 0);
    signal NK_612_583_buffered : std_logic_vector(31 downto 0);
    signal NL_730 : std_logic_vector(11 downto 0);
    signal NL_730_571_buffered : std_logic_vector(11 downto 0);
    signal NNG_478 : std_logic_vector(31 downto 0);
    signal NNJ_486 : std_logic_vector(31 downto 0);
    signal NNNT_359 : std_logic_vector(11 downto 0);
    signal NNT_369 : std_logic_vector(31 downto 0);
    signal NTT_364 : std_logic_vector(30 downto 0);
    signal NT_437 : std_logic_vector(11 downto 0);
    signal NT_437_350_buffered : std_logic_vector(11 downto 0);
    signal PJ_440_delayed_7_0_506 : std_logic_vector(15 downto 0);
    signal PPJ_444_delayed_6_0_513 : std_logic_vector(15 downto 0);
    signal PPJ_503 : std_logic_vector(15 downto 0);
    signal PPPJ_466_delayed_6_0_538 : std_logic_vector(15 downto 0);
    signal PPPJ_530 : std_logic_vector(15 downto 0);
    signal PPPPJ_470_delayed_6_0_545 : std_logic_vector(15 downto 0);
    signal PPPPJ_535 : std_logic_vector(15 downto 0);
    signal R_HHHH_684_resized : std_logic_vector(3 downto 0);
    signal R_HHHH_684_scaled : std_logic_vector(3 downto 0);
    signal R_HHH_594_delayed_4_0_682_resized : std_logic_vector(3 downto 0);
    signal R_HHH_594_delayed_4_0_682_scaled : std_logic_vector(3 downto 0);
    signal R_HHH_671_resized : std_logic_vector(3 downto 0);
    signal R_HHH_671_scaled : std_logic_vector(3 downto 0);
    signal R_HH_584_delayed_4_0_669_resized : std_logic_vector(3 downto 0);
    signal R_HH_584_delayed_4_0_669_scaled : std_logic_vector(3 downto 0);
    signal R_HH_658_resized : std_logic_vector(3 downto 0);
    signal R_HH_658_scaled : std_logic_vector(3 downto 0);
    signal R_H_574_delayed_5_0_656_resized : std_logic_vector(3 downto 0);
    signal R_H_574_delayed_5_0_656_scaled : std_logic_vector(3 downto 0);
    signal R_K_517_delayed_5_0_596_resized : std_logic_vector(3 downto 0);
    signal R_K_517_delayed_5_0_596_scaled : std_logic_vector(3 downto 0);
    signal R_K_586_resized : std_logic_vector(3 downto 0);
    signal R_K_586_scaled : std_logic_vector(3 downto 0);
    signal R_K_590_resized : std_logic_vector(3 downto 0);
    signal R_K_590_scaled : std_logic_vector(3 downto 0);
    signal R_K_604_resized : std_logic_vector(3 downto 0);
    signal R_K_604_scaled : std_logic_vector(3 downto 0);
    signal R_PJ_440_delayed_7_0_507_resized : std_logic_vector(3 downto 0);
    signal R_PJ_440_delayed_7_0_507_scaled : std_logic_vector(3 downto 0);
    signal R_PPJ_444_delayed_6_0_514_resized : std_logic_vector(3 downto 0);
    signal R_PPJ_444_delayed_6_0_514_scaled : std_logic_vector(3 downto 0);
    signal R_PPPJ_466_delayed_6_0_539_resized : std_logic_vector(3 downto 0);
    signal R_PPPJ_466_delayed_6_0_539_scaled : std_logic_vector(3 downto 0);
    signal R_PPPPJ_470_delayed_6_0_546_resized : std_logic_vector(3 downto 0);
    signal R_PPPPJ_470_delayed_6_0_546_scaled : std_logic_vector(3 downto 0);
    signal R_TTTT_371_delayed_11_0_429_resized : std_logic_vector(3 downto 0);
    signal R_TTTT_371_delayed_11_0_429_scaled : std_logic_vector(3 downto 0);
    signal R_TTT_367_delayed_11_0_422_resized : std_logic_vector(3 downto 0);
    signal R_TTT_367_delayed_11_0_422_scaled : std_logic_vector(3 downto 0);
    signal R_TT_345_delayed_11_0_397_resized : std_logic_vector(3 downto 0);
    signal R_TT_345_delayed_11_0_397_scaled : std_logic_vector(3 downto 0);
    signal R_T_341_delayed_12_0_390_resized : std_logic_vector(3 downto 0);
    signal R_T_341_delayed_12_0_390_scaled : std_logic_vector(3 downto 0);
    signal R_f_636_resized : std_logic_vector(10 downto 0);
    signal R_f_636_scaled : std_logic_vector(10 downto 0);
    signal STORE_PJ_451_data_0 : std_logic_vector(15 downto 0);
    signal STORE_PJ_451_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_PJ_555_data_0 : std_logic_vector(15 downto 0);
    signal STORE_PJ_555_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_total_573_data_0 : std_logic_vector(15 downto 0);
    signal STORE_total_573_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_total_602_data_0 : std_logic_vector(15 downto 0);
    signal STORE_total_602_word_address_0 : std_logic_vector(0 downto 0);
    signal TTTT_371_delayed_11_0_428 : std_logic_vector(11 downto 0);
    signal TTTT_418 : std_logic_vector(11 downto 0);
    signal TTT_367_delayed_11_0_421 : std_logic_vector(11 downto 0);
    signal TTT_413 : std_logic_vector(11 downto 0);
    signal TT_345_delayed_11_0_396 : std_logic_vector(11 downto 0);
    signal TT_386 : std_logic_vector(11 downto 0);
    signal T_310_delayed_4_0_354 : std_logic_vector(11 downto 0);
    signal T_341_delayed_12_0_389 : std_logic_vector(11 downto 0);
    signal T_346 : std_logic_vector(11 downto 0);
    signal ULT_u12_u1_441_wire : std_logic_vector(0 downto 0);
    signal ULT_u12_u1_563_wire : std_logic_vector(0 downto 0);
    signal ULT_u12_u1_695_wire : std_logic_vector(0 downto 0);
    signal ULT_u12_u1_734_wire : std_logic_vector(0 downto 0);
    signal ULT_u12_u1_746_wire : std_logic_vector(0 downto 0);
    signal ULT_u32_u1_616_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_391_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_391_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_391_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_391_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_391_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_391_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_391_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_398_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_398_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_398_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_398_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_398_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_398_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_398_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_423_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_423_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_423_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_423_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_423_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_423_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_423_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_430_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_430_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_430_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_430_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_430_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_430_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_430_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_508_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_508_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_508_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_508_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_508_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_508_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_508_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_515_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_515_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_515_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_515_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_515_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_515_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_515_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_540_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_540_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_540_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_540_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_540_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_540_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_540_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_547_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_547_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_547_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_547_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_547_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_547_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_547_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_587_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_587_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_587_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_587_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_587_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_587_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_587_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_591_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_591_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_591_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_591_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_591_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_591_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_591_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_597_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_597_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_597_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_597_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_597_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_597_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_597_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_605_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_605_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_605_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_605_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_605_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_605_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_605_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_605_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_637_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_637_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_637_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_637_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_637_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_637_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_637_word_address_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_637_word_offset_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_657_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_657_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_657_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_657_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_657_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_657_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_657_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_659_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_659_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_659_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_659_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_659_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_659_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_659_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_659_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_670_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_670_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_670_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_670_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_670_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_670_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_670_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_672_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_672_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_672_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_672_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_672_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_672_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_672_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_672_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_683_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_683_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_683_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_683_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_683_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_683_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_683_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_685_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_685_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_685_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_685_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_685_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_685_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_685_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_685_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_707_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_707_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_712_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_712_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_717_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_717_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_722_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_722_word_address_0 : std_logic_vector(3 downto 0);
    signal f_631 : std_logic_vector(15 downto 0);
    signal imag1_588 : std_logic_vector(15 downto 0);
    signal ker1_592 : std_logic_vector(15 downto 0);
    signal konst_384_wire_constant : std_logic_vector(11 downto 0);
    signal konst_411_wire_constant : std_logic_vector(11 downto 0);
    signal konst_416_wire_constant : std_logic_vector(11 downto 0);
    signal konst_435_wire_constant : std_logic_vector(11 downto 0);
    signal konst_440_wire_constant : std_logic_vector(11 downto 0);
    signal konst_452_wire_constant : std_logic_vector(15 downto 0);
    signal konst_501_wire_constant : std_logic_vector(15 downto 0);
    signal konst_528_wire_constant : std_logic_vector(15 downto 0);
    signal konst_533_wire_constant : std_logic_vector(15 downto 0);
    signal konst_552_wire_constant : std_logic_vector(11 downto 0);
    signal konst_557_wire_constant : std_logic_vector(15 downto 0);
    signal konst_562_wire_constant : std_logic_vector(11 downto 0);
    signal konst_574_wire_constant : std_logic_vector(15 downto 0);
    signal konst_610_wire_constant : std_logic_vector(31 downto 0);
    signal konst_615_wire_constant : std_logic_vector(31 downto 0);
    signal konst_618_wire_constant : std_logic_vector(0 downto 0);
    signal konst_650_wire_constant : std_logic_vector(11 downto 0);
    signal konst_663_wire_constant : std_logic_vector(11 downto 0);
    signal konst_676_wire_constant : std_logic_vector(11 downto 0);
    signal konst_689_wire_constant : std_logic_vector(11 downto 0);
    signal konst_694_wire_constant : std_logic_vector(11 downto 0);
    signal konst_697_wire_constant : std_logic_vector(0 downto 0);
    signal konst_701_wire_constant : std_logic_vector(11 downto 0);
    signal konst_703_wire_constant : std_logic_vector(15 downto 0);
    signal konst_728_wire_constant : std_logic_vector(11 downto 0);
    signal konst_733_wire_constant : std_logic_vector(11 downto 0);
    signal konst_740_wire_constant : std_logic_vector(11 downto 0);
    signal konst_745_wire_constant : std_logic_vector(11 downto 0);
    signal rdata_624 : std_logic_vector(63 downto 0);
    signal rdatah_490 : std_logic_vector(31 downto 0);
    signal rdatahk_373 : std_logic_vector(31 downto 0);
    signal rdatai0_498 : std_logic_vector(15 downto 0);
    signal rdatai1_494 : std_logic_vector(15 downto 0);
    signal rdatai2_525 : std_logic_vector(15 downto 0);
    signal rdatai3_521 : std_logic_vector(15 downto 0);
    signal rdatak0_381 : std_logic_vector(15 downto 0);
    signal rdatak1_377 : std_logic_vector(15 downto 0);
    signal rdatak2_408 : std_logic_vector(15 downto 0);
    signal rdatak3_404 : std_logic_vector(15 downto 0);
    signal rdatal_490 : std_logic_vector(31 downto 0);
    signal rdatalk_373 : std_logic_vector(31 downto 0);
    signal rdatar_705 : std_logic_vector(63 downto 0);
    signal slice_709_wire : std_logic_vector(15 downto 0);
    signal slice_714_wire : std_logic_vector(15 downto 0);
    signal slice_719_wire : std_logic_vector(15 downto 0);
    signal slice_724_wire : std_logic_vector(15 downto 0);
    signal type_cast_349_wire_constant : std_logic_vector(11 downto 0);
    signal type_cast_448_wire_constant : std_logic_vector(11 downto 0);
    signal type_cast_460_wire_constant : std_logic_vector(11 downto 0);
    signal type_cast_570_wire_constant : std_logic_vector(11 downto 0);
    signal type_cast_582_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_645_wire_constant : std_logic_vector(11 downto 0);
    -- 
  begin -- 
    LOAD_PJ_500_word_address_0 <= "0";
    LOAD_PJ_505_word_address_0 <= "0";
    LOAD_PJ_527_word_address_0 <= "0";
    LOAD_PJ_532_word_address_0 <= "0";
    LOAD_PJ_556_word_address_0 <= "0";
    LOAD_ZJ_357_word_address_0 <= "0";
    LOAD_one_366_word_address_0 <= "0";
    LOAD_one_475_word_address_0 <= "0";
    LOAD_total_603_word_address_0 <= "0";
    LOAD_total_622_word_address_0 <= "0";
    LOAD_zer_626_word_address_0 <= "0";
    STORE_PJ_451_word_address_0 <= "0";
    STORE_PJ_555_word_address_0 <= "0";
    STORE_total_573_word_address_0 <= "0";
    STORE_total_602_word_address_0 <= "0";
    array_obj_ref_391_offset_scale_factor_0 <= "0001";
    array_obj_ref_391_resized_base_address <= "0000";
    array_obj_ref_391_word_offset_0 <= "0000";
    array_obj_ref_398_offset_scale_factor_0 <= "0001";
    array_obj_ref_398_resized_base_address <= "0000";
    array_obj_ref_398_word_offset_0 <= "0000";
    array_obj_ref_423_offset_scale_factor_0 <= "0001";
    array_obj_ref_423_resized_base_address <= "0000";
    array_obj_ref_423_word_offset_0 <= "0000";
    array_obj_ref_430_offset_scale_factor_0 <= "0001";
    array_obj_ref_430_resized_base_address <= "0000";
    array_obj_ref_430_word_offset_0 <= "0000";
    array_obj_ref_508_offset_scale_factor_0 <= "0001";
    array_obj_ref_508_resized_base_address <= "0000";
    array_obj_ref_508_word_offset_0 <= "0000";
    array_obj_ref_515_offset_scale_factor_0 <= "0001";
    array_obj_ref_515_resized_base_address <= "0000";
    array_obj_ref_515_word_offset_0 <= "0000";
    array_obj_ref_540_offset_scale_factor_0 <= "0001";
    array_obj_ref_540_resized_base_address <= "0000";
    array_obj_ref_540_word_offset_0 <= "0000";
    array_obj_ref_547_offset_scale_factor_0 <= "0001";
    array_obj_ref_547_resized_base_address <= "0000";
    array_obj_ref_547_word_offset_0 <= "0000";
    array_obj_ref_587_offset_scale_factor_0 <= "0001";
    array_obj_ref_587_resized_base_address <= "0000";
    array_obj_ref_587_word_offset_0 <= "0000";
    array_obj_ref_591_offset_scale_factor_0 <= "0001";
    array_obj_ref_591_resized_base_address <= "0000";
    array_obj_ref_591_word_offset_0 <= "0000";
    array_obj_ref_597_offset_scale_factor_0 <= "0001";
    array_obj_ref_597_resized_base_address <= "0000";
    array_obj_ref_597_word_offset_0 <= "0000";
    array_obj_ref_605_offset_scale_factor_0 <= "0001";
    array_obj_ref_605_resized_base_address <= "0000";
    array_obj_ref_605_word_offset_0 <= "0000";
    array_obj_ref_637_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_637_resized_base_address <= "00000000000";
    array_obj_ref_637_word_offset_0 <= "00000000000";
    array_obj_ref_657_offset_scale_factor_0 <= "0001";
    array_obj_ref_657_resized_base_address <= "0000";
    array_obj_ref_657_word_offset_0 <= "0000";
    array_obj_ref_659_offset_scale_factor_0 <= "0001";
    array_obj_ref_659_resized_base_address <= "0000";
    array_obj_ref_659_word_offset_0 <= "0000";
    array_obj_ref_670_offset_scale_factor_0 <= "0001";
    array_obj_ref_670_resized_base_address <= "0000";
    array_obj_ref_670_word_offset_0 <= "0000";
    array_obj_ref_672_offset_scale_factor_0 <= "0001";
    array_obj_ref_672_resized_base_address <= "0000";
    array_obj_ref_672_word_offset_0 <= "0000";
    array_obj_ref_683_offset_scale_factor_0 <= "0001";
    array_obj_ref_683_resized_base_address <= "0000";
    array_obj_ref_683_word_offset_0 <= "0000";
    array_obj_ref_685_offset_scale_factor_0 <= "0001";
    array_obj_ref_685_resized_base_address <= "0000";
    array_obj_ref_685_word_offset_0 <= "0000";
    array_obj_ref_707_word_address_0 <= "1111";
    array_obj_ref_712_word_address_0 <= "1011";
    array_obj_ref_717_word_address_0 <= "0111";
    array_obj_ref_722_word_address_0 <= "0011";
    konst_384_wire_constant <= "000000000001";
    konst_411_wire_constant <= "000000000010";
    konst_416_wire_constant <= "000000000011";
    konst_435_wire_constant <= "000000000100";
    konst_440_wire_constant <= "000000010000";
    konst_452_wire_constant <= "0000000000000000";
    konst_501_wire_constant <= "0000000000000001";
    konst_528_wire_constant <= "0000000000000010";
    konst_533_wire_constant <= "0000000000000011";
    konst_552_wire_constant <= "000000100000";
    konst_557_wire_constant <= "0000000000000100";
    konst_562_wire_constant <= "000010000000";
    konst_574_wire_constant <= "0000000000000000";
    konst_610_wire_constant <= "00000000000000000000000000000001";
    konst_615_wire_constant <= "00000000000000000000000000010000";
    konst_618_wire_constant <= "0";
    konst_650_wire_constant <= "000000000001";
    konst_663_wire_constant <= "000000000010";
    konst_676_wire_constant <= "000000000011";
    konst_689_wire_constant <= "000000000100";
    konst_694_wire_constant <= "000000010000";
    konst_697_wire_constant <= "1";
    konst_701_wire_constant <= "000000000100";
    konst_703_wire_constant <= "0000000000000000";
    konst_728_wire_constant <= "000000000001";
    konst_733_wire_constant <= "000000011101";
    konst_740_wire_constant <= "000000100000";
    konst_745_wire_constant <= "001110100000";
    type_cast_349_wire_constant <= "000000000000";
    type_cast_448_wire_constant <= "000000000000";
    type_cast_460_wire_constant <= "000000000000";
    type_cast_570_wire_constant <= "000000000000";
    type_cast_582_wire_constant <= "00000000000000000000000000000000";
    type_cast_645_wire_constant <= "000000000000";
    -- logger for phi phi_stmt_346
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_346_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:try1:DP:phi_stmt_346:input-0 type_cast_349_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_349_wire_constant));
          --
        end if;
        if phi_stmt_346_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:try1:DP:phi_stmt_346:input-1 NT_437_350_buffered= " & Convert_SLV_To_Hex_String(NT_437_350_buffered));
          --
        end if;
        if phi_stmt_346_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:try1:DP:phi_stmt_346:sample-completed");
          --
        end if;
        if phi_stmt_346_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:try1:DP:phi_stmt_346:output T_346= " & Convert_SLV_To_Hex_String(T_346));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_346: Block -- phi operator 
      signal idata: std_logic_vector(23 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_349_wire_constant & NT_437_350_buffered;
      req <= phi_stmt_346_req_0 & phi_stmt_346_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_346",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 12) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_346_ack_0,
          idata => idata,
          odata => T_346,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_346
    -- logger for phi phi_stmt_445
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_445_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:try1:DP:phi_stmt_445:input-0 type_cast_448_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_448_wire_constant));
          --
        end if;
        if phi_stmt_445_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:try1:DP:phi_stmt_445:input-1 NG_742_449_buffered= " & Convert_SLV_To_Hex_String(NG_742_449_buffered));
          --
        end if;
        if phi_stmt_445_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:try1:DP:phi_stmt_445:sample-completed");
          --
        end if;
        if phi_stmt_445_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:try1:DP:phi_stmt_445:output G_445= " & Convert_SLV_To_Hex_String(G_445));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_445: Block -- phi operator 
      signal idata: std_logic_vector(23 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_448_wire_constant & NG_742_449_buffered;
      req <= phi_stmt_445_req_0 & phi_stmt_445_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_445",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 12) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_445_ack_0,
          idata => idata,
          odata => G_445,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_445
    -- logger for phi phi_stmt_457
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_457_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:try1:DP:phi_stmt_457:input-0 type_cast_460_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_460_wire_constant));
          --
        end if;
        if phi_stmt_457_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:try1:DP:phi_stmt_457:input-1 NJ_554_461_buffered= " & Convert_SLV_To_Hex_String(NJ_554_461_buffered));
          --
        end if;
        if phi_stmt_457_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:try1:DP:phi_stmt_457:sample-completed");
          --
        end if;
        if phi_stmt_457_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:try1:DP:phi_stmt_457:output J_457= " & Convert_SLV_To_Hex_String(J_457));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_457: Block -- phi operator 
      signal idata: std_logic_vector(23 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_460_wire_constant & NJ_554_461_buffered;
      req <= phi_stmt_457_req_0 & phi_stmt_457_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_457",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 12) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_457_ack_0,
          idata => idata,
          odata => J_457,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_457
    -- logger for phi phi_stmt_567
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_567_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:try1:DP:phi_stmt_567:input-0 type_cast_570_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_570_wire_constant));
          --
        end if;
        if phi_stmt_567_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:try1:DP:phi_stmt_567:input-1 NL_730_571_buffered= " & Convert_SLV_To_Hex_String(NL_730_571_buffered));
          --
        end if;
        if phi_stmt_567_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:try1:DP:phi_stmt_567:sample-completed");
          --
        end if;
        if phi_stmt_567_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:try1:DP:phi_stmt_567:output L_567= " & Convert_SLV_To_Hex_String(L_567));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_567: Block -- phi operator 
      signal idata: std_logic_vector(23 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_570_wire_constant & NL_730_571_buffered;
      req <= phi_stmt_567_req_0 & phi_stmt_567_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_567",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 12) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_567_ack_0,
          idata => idata,
          odata => L_567,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_567
    -- logger for phi phi_stmt_579
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_579_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:try1:DP:phi_stmt_579:input-0 type_cast_582_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_582_wire_constant));
          --
        end if;
        if phi_stmt_579_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:try1:DP:phi_stmt_579:input-1 NK_612_583_buffered= " & Convert_SLV_To_Hex_String(NK_612_583_buffered));
          --
        end if;
        if phi_stmt_579_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:try1:DP:phi_stmt_579:sample-completed");
          --
        end if;
        if phi_stmt_579_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:try1:DP:phi_stmt_579:output K_579= " & Convert_SLV_To_Hex_String(K_579));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_579: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_582_wire_constant & NK_612_583_buffered;
      req <= phi_stmt_579_req_0 & phi_stmt_579_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_579",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_579_ack_0,
          idata => idata,
          odata => K_579,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_579
    -- logger for phi phi_stmt_642
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_642_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:try1:DP:phi_stmt_642:input-0 type_cast_645_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_645_wire_constant));
          --
        end if;
        if phi_stmt_642_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:try1:DP:phi_stmt_642:input-1 NH_691_646_buffered= " & Convert_SLV_To_Hex_String(NH_691_646_buffered));
          --
        end if;
        if phi_stmt_642_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:try1:DP:phi_stmt_642:sample-completed");
          --
        end if;
        if phi_stmt_642_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:try1:DP:phi_stmt_642:output H_642= " & Convert_SLV_To_Hex_String(H_642));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_642: Block -- phi operator 
      signal idata: std_logic_vector(23 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_645_wire_constant & NH_691_646_buffered;
      req <= phi_stmt_642_req_0 & phi_stmt_642_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_642",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 12) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_642_ack_0,
          idata => idata,
          odata => H_642,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_642
    -- logger for split-operator slice_376_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_376_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_376_inst:started:   inputs: " & " rdatalk_373 = "& Convert_SLV_To_Hex_String(rdatalk_373));
          --
        end if; 
        if slice_376_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_376_inst:finished:  outputs: " & " rdatak1_377= "  & Convert_SLV_To_Hex_String(rdatak1_377));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_376_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_376_inst_req_0;
      slice_376_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_376_inst_req_1;
      slice_376_inst_ack_1<= update_ack(0);
      slice_376_inst: SliceSplitProtocol generic map(name => "slice_376_inst", in_data_width => 32, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => rdatalk_373, dout => rdatak1_377, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_380_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_380_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_380_inst:started:   inputs: " & " rdatalk_373 = "& Convert_SLV_To_Hex_String(rdatalk_373));
          --
        end if; 
        if slice_380_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_380_inst:finished:  outputs: " & " rdatak0_381= "  & Convert_SLV_To_Hex_String(rdatak0_381));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_380_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_380_inst_req_0;
      slice_380_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_380_inst_req_1;
      slice_380_inst_ack_1<= update_ack(0);
      slice_380_inst: SliceSplitProtocol generic map(name => "slice_380_inst", in_data_width => 32, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => rdatalk_373, dout => rdatak0_381, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_403_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_403_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_403_inst:started:   inputs: " & " rdatahk_373 = "& Convert_SLV_To_Hex_String(rdatahk_373));
          --
        end if; 
        if slice_403_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_403_inst:finished:  outputs: " & " rdatak3_404= "  & Convert_SLV_To_Hex_String(rdatak3_404));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_403_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_403_inst_req_0;
      slice_403_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_403_inst_req_1;
      slice_403_inst_ack_1<= update_ack(0);
      slice_403_inst: SliceSplitProtocol generic map(name => "slice_403_inst", in_data_width => 32, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => rdatahk_373, dout => rdatak3_404, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_407_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_407_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_407_inst:started:   inputs: " & " rdatahk_373 = "& Convert_SLV_To_Hex_String(rdatahk_373));
          --
        end if; 
        if slice_407_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_407_inst:finished:  outputs: " & " rdatak2_408= "  & Convert_SLV_To_Hex_String(rdatak2_408));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_407_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_407_inst_req_0;
      slice_407_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_407_inst_req_1;
      slice_407_inst_ack_1<= update_ack(0);
      slice_407_inst: SliceSplitProtocol generic map(name => "slice_407_inst", in_data_width => 32, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => rdatahk_373, dout => rdatak2_408, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_493_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_493_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_493_inst:started:   inputs: " & " rdatal_490 = "& Convert_SLV_To_Hex_String(rdatal_490));
          --
        end if; 
        if slice_493_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_493_inst:finished:  outputs: " & " rdatai1_494= "  & Convert_SLV_To_Hex_String(rdatai1_494));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_493_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_493_inst_req_0;
      slice_493_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_493_inst_req_1;
      slice_493_inst_ack_1<= update_ack(0);
      slice_493_inst: SliceSplitProtocol generic map(name => "slice_493_inst", in_data_width => 32, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => rdatal_490, dout => rdatai1_494, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_497_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_497_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_497_inst:started:   inputs: " & " rdatal_490 = "& Convert_SLV_To_Hex_String(rdatal_490));
          --
        end if; 
        if slice_497_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_497_inst:finished:  outputs: " & " rdatai0_498= "  & Convert_SLV_To_Hex_String(rdatai0_498));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_497_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_497_inst_req_0;
      slice_497_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_497_inst_req_1;
      slice_497_inst_ack_1<= update_ack(0);
      slice_497_inst: SliceSplitProtocol generic map(name => "slice_497_inst", in_data_width => 32, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => rdatal_490, dout => rdatai0_498, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_520_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_520_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_520_inst:started:   inputs: " & " rdatah_490 = "& Convert_SLV_To_Hex_String(rdatah_490));
          --
        end if; 
        if slice_520_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_520_inst:finished:  outputs: " & " rdatai3_521= "  & Convert_SLV_To_Hex_String(rdatai3_521));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_520_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_520_inst_req_0;
      slice_520_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_520_inst_req_1;
      slice_520_inst_ack_1<= update_ack(0);
      slice_520_inst: SliceSplitProtocol generic map(name => "slice_520_inst", in_data_width => 32, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => rdatah_490, dout => rdatai3_521, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_524_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_524_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_524_inst:started:   inputs: " & " rdatah_490 = "& Convert_SLV_To_Hex_String(rdatah_490));
          --
        end if; 
        if slice_524_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_524_inst:finished:  outputs: " & " rdatai2_525= "  & Convert_SLV_To_Hex_String(rdatai2_525));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_524_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_524_inst_req_0;
      slice_524_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_524_inst_req_1;
      slice_524_inst_ack_1<= update_ack(0);
      slice_524_inst: SliceSplitProtocol generic map(name => "slice_524_inst", in_data_width => 32, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => rdatah_490, dout => rdatai2_525, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_709_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_709_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_709_inst:started:   inputs: " & " rdatar_705 = "& Convert_SLV_To_Hex_String(rdatar_705));
          --
        end if; 
        if slice_709_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_709_inst:finished:  outputs: " & " slice_709_wire= "  & Convert_SLV_To_Hex_String(slice_709_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_709_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_709_inst_req_0;
      slice_709_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_709_inst_req_1;
      slice_709_inst_ack_1<= update_ack(0);
      slice_709_inst: SliceSplitProtocol generic map(name => "slice_709_inst", in_data_width => 64, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => rdatar_705, dout => slice_709_wire, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_714_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_714_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_714_inst:started:   inputs: " & " rdatar_705 = "& Convert_SLV_To_Hex_String(rdatar_705));
          --
        end if; 
        if slice_714_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_714_inst:finished:  outputs: " & " slice_714_wire= "  & Convert_SLV_To_Hex_String(slice_714_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_714_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_714_inst_req_0;
      slice_714_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_714_inst_req_1;
      slice_714_inst_ack_1<= update_ack(0);
      slice_714_inst: SliceSplitProtocol generic map(name => "slice_714_inst", in_data_width => 64, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => rdatar_705, dout => slice_714_wire, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_719_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_719_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_719_inst:started:   inputs: " & " rdatar_705 = "& Convert_SLV_To_Hex_String(rdatar_705));
          --
        end if; 
        if slice_719_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_719_inst:finished:  outputs: " & " slice_719_wire= "  & Convert_SLV_To_Hex_String(slice_719_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_719_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_719_inst_req_0;
      slice_719_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_719_inst_req_1;
      slice_719_inst_ack_1<= update_ack(0);
      slice_719_inst: SliceSplitProtocol generic map(name => "slice_719_inst", in_data_width => 64, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => rdatar_705, dout => slice_719_wire, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_724_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_724_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_724_inst:started:   inputs: " & " rdatar_705 = "& Convert_SLV_To_Hex_String(rdatar_705));
          --
        end if; 
        if slice_724_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:slice_724_inst:finished:  outputs: " & " slice_724_wire= "  & Convert_SLV_To_Hex_String(slice_724_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_724_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_724_inst_req_0;
      slice_724_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_724_inst_req_1;
      slice_724_inst_ack_1<= update_ack(0);
      slice_724_inst: SliceSplitProtocol generic map(name => "slice_724_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => rdatar_705, dout => slice_724_wire, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator NG_742_449_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if NG_742_449_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:NG_742_449_buf:started:   inputs: " & " NG_742 = "& Convert_SLV_To_Hex_String(NG_742));
          --
        end if; 
        if NG_742_449_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:NG_742_449_buf:finished:  outputs: " & " NG_742_449_buffered= "  & Convert_SLV_To_Hex_String(NG_742_449_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    NG_742_449_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= NG_742_449_buf_req_0;
      NG_742_449_buf_ack_0<= wack(0);
      rreq(0) <= NG_742_449_buf_req_1;
      NG_742_449_buf_ack_1<= rack(0);
      NG_742_449_buf : InterlockBuffer generic map ( -- 
        name => "NG_742_449_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => NG_742,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NG_742_449_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator NH_691_646_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if NH_691_646_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:NH_691_646_buf:started:   inputs: " & " NH_691 = "& Convert_SLV_To_Hex_String(NH_691));
          --
        end if; 
        if NH_691_646_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:NH_691_646_buf:finished:  outputs: " & " NH_691_646_buffered= "  & Convert_SLV_To_Hex_String(NH_691_646_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    NH_691_646_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= NH_691_646_buf_req_0;
      NH_691_646_buf_ack_0<= wack(0);
      rreq(0) <= NH_691_646_buf_req_1;
      NH_691_646_buf_ack_1<= rack(0);
      NH_691_646_buf : InterlockBuffer generic map ( -- 
        name => "NH_691_646_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => NH_691,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NH_691_646_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator NJ_554_461_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if NJ_554_461_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:NJ_554_461_buf:started:   inputs: " & " NJ_554 = "& Convert_SLV_To_Hex_String(NJ_554));
          --
        end if; 
        if NJ_554_461_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:NJ_554_461_buf:finished:  outputs: " & " NJ_554_461_buffered= "  & Convert_SLV_To_Hex_String(NJ_554_461_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    NJ_554_461_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= NJ_554_461_buf_req_0;
      NJ_554_461_buf_ack_0<= wack(0);
      rreq(0) <= NJ_554_461_buf_req_1;
      NJ_554_461_buf_ack_1<= rack(0);
      NJ_554_461_buf : InterlockBuffer generic map ( -- 
        name => "NJ_554_461_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => NJ_554,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NJ_554_461_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator NK_612_583_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if NK_612_583_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:NK_612_583_buf:started:   inputs: " & " NK_612 = "& Convert_SLV_To_Hex_String(NK_612));
          --
        end if; 
        if NK_612_583_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:NK_612_583_buf:finished:  outputs: " & " NK_612_583_buffered= "  & Convert_SLV_To_Hex_String(NK_612_583_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    NK_612_583_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= NK_612_583_buf_req_0;
      NK_612_583_buf_ack_0<= wack(0);
      rreq(0) <= NK_612_583_buf_req_1;
      NK_612_583_buf_ack_1<= rack(0);
      NK_612_583_buf : InterlockBuffer generic map ( -- 
        name => "NK_612_583_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => NK_612,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NK_612_583_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator NL_730_571_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if NL_730_571_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:NL_730_571_buf:started:   inputs: " & " NL_730 = "& Convert_SLV_To_Hex_String(NL_730));
          --
        end if; 
        if NL_730_571_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:NL_730_571_buf:finished:  outputs: " & " NL_730_571_buffered= "  & Convert_SLV_To_Hex_String(NL_730_571_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    NL_730_571_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= NL_730_571_buf_req_0;
      NL_730_571_buf_ack_0<= wack(0);
      rreq(0) <= NL_730_571_buf_req_1;
      NL_730_571_buf_ack_1<= rack(0);
      NL_730_571_buf : InterlockBuffer generic map ( -- 
        name => "NL_730_571_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => NL_730,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NL_730_571_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator NT_437_350_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if NT_437_350_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:NT_437_350_buf:started:   inputs: " & " NT_437 = "& Convert_SLV_To_Hex_String(NT_437));
          --
        end if; 
        if NT_437_350_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:NT_437_350_buf:finished:  outputs: " & " NT_437_350_buffered= "  & Convert_SLV_To_Hex_String(NT_437_350_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    NT_437_350_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= NT_437_350_buf_req_0;
      NT_437_350_buf_ack_0<= wack(0);
      rreq(0) <= NT_437_350_buf_req_1;
      NT_437_350_buf_ack_1<= rack(0);
      NT_437_350_buf : InterlockBuffer generic map ( -- 
        name => "NT_437_350_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => NT_437,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NT_437_350_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_HHH_594_delayed_4_0_679_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_HHH_594_delayed_4_0_679_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_HHH_594_delayed_4_0_679_inst:started:   inputs: " & " HHH_665 = "& Convert_SLV_To_Hex_String(HHH_665));
          --
        end if; 
        if W_HHH_594_delayed_4_0_679_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_HHH_594_delayed_4_0_679_inst:finished:  outputs: " & " HHH_594_delayed_4_0_681= "  & Convert_SLV_To_Hex_String(HHH_594_delayed_4_0_681));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_HHH_594_delayed_4_0_679_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_HHH_594_delayed_4_0_679_inst_req_0;
      W_HHH_594_delayed_4_0_679_inst_ack_0<= wack(0);
      rreq(0) <= W_HHH_594_delayed_4_0_679_inst_req_1;
      W_HHH_594_delayed_4_0_679_inst_ack_1<= rack(0);
      W_HHH_594_delayed_4_0_679_inst : InterlockBuffer generic map ( -- 
        name => "W_HHH_594_delayed_4_0_679_inst",
        buffer_size => 4,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => HHH_665,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => HHH_594_delayed_4_0_681,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_HH_584_delayed_4_0_666_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_HH_584_delayed_4_0_666_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_HH_584_delayed_4_0_666_inst:started:   inputs: " & " HH_652 = "& Convert_SLV_To_Hex_String(HH_652));
          --
        end if; 
        if W_HH_584_delayed_4_0_666_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_HH_584_delayed_4_0_666_inst:finished:  outputs: " & " HH_584_delayed_4_0_668= "  & Convert_SLV_To_Hex_String(HH_584_delayed_4_0_668));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_HH_584_delayed_4_0_666_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_HH_584_delayed_4_0_666_inst_req_0;
      W_HH_584_delayed_4_0_666_inst_ack_0<= wack(0);
      rreq(0) <= W_HH_584_delayed_4_0_666_inst_req_1;
      W_HH_584_delayed_4_0_666_inst_ack_1<= rack(0);
      W_HH_584_delayed_4_0_666_inst : InterlockBuffer generic map ( -- 
        name => "W_HH_584_delayed_4_0_666_inst",
        buffer_size => 4,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => HH_652,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => HH_584_delayed_4_0_668,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_H_574_delayed_5_0_653_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_H_574_delayed_5_0_653_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_H_574_delayed_5_0_653_inst:started:   inputs: " & " H_642 = "& Convert_SLV_To_Hex_String(H_642));
          --
        end if; 
        if W_H_574_delayed_5_0_653_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_H_574_delayed_5_0_653_inst:finished:  outputs: " & " H_574_delayed_5_0_655= "  & Convert_SLV_To_Hex_String(H_574_delayed_5_0_655));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_H_574_delayed_5_0_653_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_H_574_delayed_5_0_653_inst_req_0;
      W_H_574_delayed_5_0_653_inst_ack_0<= wack(0);
      rreq(0) <= W_H_574_delayed_5_0_653_inst_req_1;
      W_H_574_delayed_5_0_653_inst_ack_1<= rack(0);
      W_H_574_delayed_5_0_653_inst : InterlockBuffer generic map ( -- 
        name => "W_H_574_delayed_5_0_653_inst",
        buffer_size => 5,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => H_642,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => H_574_delayed_5_0_655,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_K_517_delayed_5_0_593_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_K_517_delayed_5_0_593_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_K_517_delayed_5_0_593_inst:started:   inputs: " & " K_579 = "& Convert_SLV_To_Hex_String(K_579));
          --
        end if; 
        if W_K_517_delayed_5_0_593_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_K_517_delayed_5_0_593_inst:finished:  outputs: " & " K_517_delayed_5_0_595= "  & Convert_SLV_To_Hex_String(K_517_delayed_5_0_595));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_K_517_delayed_5_0_593_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_K_517_delayed_5_0_593_inst_req_0;
      W_K_517_delayed_5_0_593_inst_ack_0<= wack(0);
      rreq(0) <= W_K_517_delayed_5_0_593_inst_req_1;
      W_K_517_delayed_5_0_593_inst_ack_1<= rack(0);
      W_K_517_delayed_5_0_593_inst : InterlockBuffer generic map ( -- 
        name => "W_K_517_delayed_5_0_593_inst",
        buffer_size => 5,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => K_579,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => K_517_delayed_5_0_595,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_NGG_420_delayed_4_0_479_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_NGG_420_delayed_4_0_479_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_NGG_420_delayed_4_0_479_inst:started:   inputs: " & " NGG_470 = "& Convert_SLV_To_Hex_String(NGG_470));
          --
        end if; 
        if W_NGG_420_delayed_4_0_479_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_NGG_420_delayed_4_0_479_inst:finished:  outputs: " & " NGG_420_delayed_4_0_481= "  & Convert_SLV_To_Hex_String(NGG_420_delayed_4_0_481));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_NGG_420_delayed_4_0_479_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_NGG_420_delayed_4_0_479_inst_req_0;
      W_NGG_420_delayed_4_0_479_inst_ack_0<= wack(0);
      rreq(0) <= W_NGG_420_delayed_4_0_479_inst_req_1;
      W_NGG_420_delayed_4_0_479_inst_ack_1<= rack(0);
      W_NGG_420_delayed_4_0_479_inst : InterlockBuffer generic map ( -- 
        name => "W_NGG_420_delayed_4_0_479_inst",
        buffer_size => 4,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => NGG_470,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NGG_420_delayed_4_0_481,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_NJJ_415_delayed_2_0_471_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_NJJ_415_delayed_2_0_471_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_NJJ_415_delayed_2_0_471_inst:started:   inputs: " & " NJJ_466 = "& Convert_SLV_To_Hex_String(NJJ_466));
          --
        end if; 
        if W_NJJ_415_delayed_2_0_471_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_NJJ_415_delayed_2_0_471_inst:finished:  outputs: " & " NJJ_415_delayed_2_0_473= "  & Convert_SLV_To_Hex_String(NJJ_415_delayed_2_0_473));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_NJJ_415_delayed_2_0_471_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_NJJ_415_delayed_2_0_471_inst_req_0;
      W_NJJ_415_delayed_2_0_471_inst_ack_0<= wack(0);
      rreq(0) <= W_NJJ_415_delayed_2_0_471_inst_req_1;
      W_NJJ_415_delayed_2_0_471_inst_ack_1<= rack(0);
      W_NJJ_415_delayed_2_0_471_inst : InterlockBuffer generic map ( -- 
        name => "W_NJJ_415_delayed_2_0_471_inst",
        buffer_size => 2,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 31,
        out_data_width => 31,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => NJJ_466,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NJJ_415_delayed_2_0_473,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_PPJ_444_delayed_6_0_511_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_PPJ_444_delayed_6_0_511_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_PPJ_444_delayed_6_0_511_inst:started:   inputs: " & " PPJ_503 = "& Convert_SLV_To_Hex_String(PPJ_503));
          --
        end if; 
        if W_PPJ_444_delayed_6_0_511_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_PPJ_444_delayed_6_0_511_inst:finished:  outputs: " & " PPJ_444_delayed_6_0_513= "  & Convert_SLV_To_Hex_String(PPJ_444_delayed_6_0_513));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_PPJ_444_delayed_6_0_511_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_PPJ_444_delayed_6_0_511_inst_req_0;
      W_PPJ_444_delayed_6_0_511_inst_ack_0<= wack(0);
      rreq(0) <= W_PPJ_444_delayed_6_0_511_inst_req_1;
      W_PPJ_444_delayed_6_0_511_inst_ack_1<= rack(0);
      W_PPJ_444_delayed_6_0_511_inst : InterlockBuffer generic map ( -- 
        name => "W_PPJ_444_delayed_6_0_511_inst",
        buffer_size => 6,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => PPJ_503,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => PPJ_444_delayed_6_0_513,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_PPPJ_466_delayed_6_0_536_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_PPPJ_466_delayed_6_0_536_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_PPPJ_466_delayed_6_0_536_inst:started:   inputs: " & " PPPJ_530 = "& Convert_SLV_To_Hex_String(PPPJ_530));
          --
        end if; 
        if W_PPPJ_466_delayed_6_0_536_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_PPPJ_466_delayed_6_0_536_inst:finished:  outputs: " & " PPPJ_466_delayed_6_0_538= "  & Convert_SLV_To_Hex_String(PPPJ_466_delayed_6_0_538));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_PPPJ_466_delayed_6_0_536_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_PPPJ_466_delayed_6_0_536_inst_req_0;
      W_PPPJ_466_delayed_6_0_536_inst_ack_0<= wack(0);
      rreq(0) <= W_PPPJ_466_delayed_6_0_536_inst_req_1;
      W_PPPJ_466_delayed_6_0_536_inst_ack_1<= rack(0);
      W_PPPJ_466_delayed_6_0_536_inst : InterlockBuffer generic map ( -- 
        name => "W_PPPJ_466_delayed_6_0_536_inst",
        buffer_size => 6,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => PPPJ_530,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => PPPJ_466_delayed_6_0_538,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_PPPPJ_470_delayed_6_0_543_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_PPPPJ_470_delayed_6_0_543_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_PPPPJ_470_delayed_6_0_543_inst:started:   inputs: " & " PPPPJ_535 = "& Convert_SLV_To_Hex_String(PPPPJ_535));
          --
        end if; 
        if W_PPPPJ_470_delayed_6_0_543_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_PPPPJ_470_delayed_6_0_543_inst:finished:  outputs: " & " PPPPJ_470_delayed_6_0_545= "  & Convert_SLV_To_Hex_String(PPPPJ_470_delayed_6_0_545));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_PPPPJ_470_delayed_6_0_543_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_PPPPJ_470_delayed_6_0_543_inst_req_0;
      W_PPPPJ_470_delayed_6_0_543_inst_ack_0<= wack(0);
      rreq(0) <= W_PPPPJ_470_delayed_6_0_543_inst_req_1;
      W_PPPPJ_470_delayed_6_0_543_inst_ack_1<= rack(0);
      W_PPPPJ_470_delayed_6_0_543_inst : InterlockBuffer generic map ( -- 
        name => "W_PPPPJ_470_delayed_6_0_543_inst",
        buffer_size => 6,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => PPPPJ_535,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => PPPPJ_470_delayed_6_0_545,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_TTTT_371_delayed_11_0_426_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_TTTT_371_delayed_11_0_426_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_TTTT_371_delayed_11_0_426_inst:started:   inputs: " & " TTTT_418 = "& Convert_SLV_To_Hex_String(TTTT_418));
          --
        end if; 
        if W_TTTT_371_delayed_11_0_426_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_TTTT_371_delayed_11_0_426_inst:finished:  outputs: " & " TTTT_371_delayed_11_0_428= "  & Convert_SLV_To_Hex_String(TTTT_371_delayed_11_0_428));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_TTTT_371_delayed_11_0_426_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_TTTT_371_delayed_11_0_426_inst_req_0;
      W_TTTT_371_delayed_11_0_426_inst_ack_0<= wack(0);
      rreq(0) <= W_TTTT_371_delayed_11_0_426_inst_req_1;
      W_TTTT_371_delayed_11_0_426_inst_ack_1<= rack(0);
      W_TTTT_371_delayed_11_0_426_inst : InterlockBuffer generic map ( -- 
        name => "W_TTTT_371_delayed_11_0_426_inst",
        buffer_size => 11,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => TTTT_418,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => TTTT_371_delayed_11_0_428,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_TTT_367_delayed_11_0_419_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_TTT_367_delayed_11_0_419_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_TTT_367_delayed_11_0_419_inst:started:   inputs: " & " TTT_413 = "& Convert_SLV_To_Hex_String(TTT_413));
          --
        end if; 
        if W_TTT_367_delayed_11_0_419_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_TTT_367_delayed_11_0_419_inst:finished:  outputs: " & " TTT_367_delayed_11_0_421= "  & Convert_SLV_To_Hex_String(TTT_367_delayed_11_0_421));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_TTT_367_delayed_11_0_419_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_TTT_367_delayed_11_0_419_inst_req_0;
      W_TTT_367_delayed_11_0_419_inst_ack_0<= wack(0);
      rreq(0) <= W_TTT_367_delayed_11_0_419_inst_req_1;
      W_TTT_367_delayed_11_0_419_inst_ack_1<= rack(0);
      W_TTT_367_delayed_11_0_419_inst : InterlockBuffer generic map ( -- 
        name => "W_TTT_367_delayed_11_0_419_inst",
        buffer_size => 11,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => TTT_413,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => TTT_367_delayed_11_0_421,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_TT_345_delayed_11_0_394_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_TT_345_delayed_11_0_394_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_TT_345_delayed_11_0_394_inst:started:   inputs: " & " TT_386 = "& Convert_SLV_To_Hex_String(TT_386));
          --
        end if; 
        if W_TT_345_delayed_11_0_394_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_TT_345_delayed_11_0_394_inst:finished:  outputs: " & " TT_345_delayed_11_0_396= "  & Convert_SLV_To_Hex_String(TT_345_delayed_11_0_396));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_TT_345_delayed_11_0_394_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_TT_345_delayed_11_0_394_inst_req_0;
      W_TT_345_delayed_11_0_394_inst_ack_0<= wack(0);
      rreq(0) <= W_TT_345_delayed_11_0_394_inst_req_1;
      W_TT_345_delayed_11_0_394_inst_ack_1<= rack(0);
      W_TT_345_delayed_11_0_394_inst : InterlockBuffer generic map ( -- 
        name => "W_TT_345_delayed_11_0_394_inst",
        buffer_size => 11,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => TT_386,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => TT_345_delayed_11_0_396,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_T_310_delayed_4_0_352_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_T_310_delayed_4_0_352_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_T_310_delayed_4_0_352_inst:started:   inputs: " & " T_346 = "& Convert_SLV_To_Hex_String(T_346));
          --
        end if; 
        if W_T_310_delayed_4_0_352_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_T_310_delayed_4_0_352_inst:finished:  outputs: " & " T_310_delayed_4_0_354= "  & Convert_SLV_To_Hex_String(T_310_delayed_4_0_354));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_T_310_delayed_4_0_352_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_T_310_delayed_4_0_352_inst_req_0;
      W_T_310_delayed_4_0_352_inst_ack_0<= wack(0);
      rreq(0) <= W_T_310_delayed_4_0_352_inst_req_1;
      W_T_310_delayed_4_0_352_inst_ack_1<= rack(0);
      W_T_310_delayed_4_0_352_inst : InterlockBuffer generic map ( -- 
        name => "W_T_310_delayed_4_0_352_inst",
        buffer_size => 4,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => T_346,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => T_310_delayed_4_0_354,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_T_341_delayed_12_0_387_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_T_341_delayed_12_0_387_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_T_341_delayed_12_0_387_inst:started:   inputs: " & " T_346 = "& Convert_SLV_To_Hex_String(T_346));
          --
        end if; 
        if W_T_341_delayed_12_0_387_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:W_T_341_delayed_12_0_387_inst:finished:  outputs: " & " T_341_delayed_12_0_389= "  & Convert_SLV_To_Hex_String(T_341_delayed_12_0_389));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_T_341_delayed_12_0_387_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_T_341_delayed_12_0_387_inst_req_0;
      W_T_341_delayed_12_0_387_inst_ack_0<= wack(0);
      rreq(0) <= W_T_341_delayed_12_0_387_inst_req_1;
      W_T_341_delayed_12_0_387_inst_ack_1<= rack(0);
      W_T_341_delayed_12_0_387_inst : InterlockBuffer generic map ( -- 
        name => "W_T_341_delayed_12_0_387_inst",
        buffer_size => 12,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => T_346,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => T_341_delayed_12_0_389,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_363_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_363_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:type_cast_363_inst:started:   inputs: " & " NNNT_359 = "& Convert_SLV_To_Hex_String(NNNT_359));
          --
        end if; 
        if type_cast_363_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:type_cast_363_inst:finished:  outputs: " & " NTT_364= "  & Convert_SLV_To_Hex_String(NTT_364));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_363_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_363_inst_req_0;
      type_cast_363_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_363_inst_req_1;
      type_cast_363_inst_ack_1<= rack(0);
      type_cast_363_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_363_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 12,
        out_data_width => 31,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => NNNT_359,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NTT_364,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_465_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_465_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:type_cast_465_inst:started:   inputs: " & " J_457 = "& Convert_SLV_To_Hex_String(J_457));
          --
        end if; 
        if type_cast_465_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:type_cast_465_inst:finished:  outputs: " & " NJJ_466= "  & Convert_SLV_To_Hex_String(NJJ_466));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_465_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_465_inst_req_0;
      type_cast_465_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_465_inst_req_1;
      type_cast_465_inst_ack_1<= rack(0);
      type_cast_465_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_465_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 12,
        out_data_width => 31,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => J_457,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NJJ_466,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_469_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_469_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:type_cast_469_inst:started:   inputs: " & " G_445 = "& Convert_SLV_To_Hex_String(G_445));
          --
        end if; 
        if type_cast_469_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:type_cast_469_inst:finished:  outputs: " & " NGG_470= "  & Convert_SLV_To_Hex_String(NGG_470));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_469_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_469_inst_req_0;
      type_cast_469_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_469_inst_req_1;
      type_cast_469_inst_ack_1<= rack(0);
      type_cast_469_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_469_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 12,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => G_445,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NGG_470,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for operator LOAD_PJ_500_gather_scatter flow-through 
    process(LOAD_PJ_500_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_PJ_500_gather_scatter:flowthrough  inputs: " & " LOAD_PJ_500_data_0 = "& Convert_SLV_To_Hex_String(LOAD_PJ_500_data_0) & "outputs: " & " LOAD_PJ_500_wire= "  & Convert_SLV_To_Hex_String(LOAD_PJ_500_wire));
      --
    end process; 
    -- equivalence LOAD_PJ_500_gather_scatter
    process(LOAD_PJ_500_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_PJ_500_data_0;
      ov(15 downto 0) := iv;
      LOAD_PJ_500_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator LOAD_PJ_505_gather_scatter flow-through 
    process(PJ_440_delayed_7_0_506) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_PJ_505_gather_scatter:flowthrough  inputs: " & " LOAD_PJ_505_data_0 = "& Convert_SLV_To_Hex_String(LOAD_PJ_505_data_0) & "outputs: " & " PJ_440_delayed_7_0_506= "  & Convert_SLV_To_Hex_String(PJ_440_delayed_7_0_506));
      --
    end process; 
    -- equivalence LOAD_PJ_505_gather_scatter
    process(LOAD_PJ_505_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_PJ_505_data_0;
      ov(15 downto 0) := iv;
      PJ_440_delayed_7_0_506 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator LOAD_PJ_527_gather_scatter flow-through 
    process(LOAD_PJ_527_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_PJ_527_gather_scatter:flowthrough  inputs: " & " LOAD_PJ_527_data_0 = "& Convert_SLV_To_Hex_String(LOAD_PJ_527_data_0) & "outputs: " & " LOAD_PJ_527_wire= "  & Convert_SLV_To_Hex_String(LOAD_PJ_527_wire));
      --
    end process; 
    -- equivalence LOAD_PJ_527_gather_scatter
    process(LOAD_PJ_527_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_PJ_527_data_0;
      ov(15 downto 0) := iv;
      LOAD_PJ_527_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator LOAD_PJ_532_gather_scatter flow-through 
    process(LOAD_PJ_532_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_PJ_532_gather_scatter:flowthrough  inputs: " & " LOAD_PJ_532_data_0 = "& Convert_SLV_To_Hex_String(LOAD_PJ_532_data_0) & "outputs: " & " LOAD_PJ_532_wire= "  & Convert_SLV_To_Hex_String(LOAD_PJ_532_wire));
      --
    end process; 
    -- equivalence LOAD_PJ_532_gather_scatter
    process(LOAD_PJ_532_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_PJ_532_data_0;
      ov(15 downto 0) := iv;
      LOAD_PJ_532_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator LOAD_PJ_556_gather_scatter flow-through 
    process(LOAD_PJ_556_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_PJ_556_gather_scatter:flowthrough  inputs: " & " LOAD_PJ_556_data_0 = "& Convert_SLV_To_Hex_String(LOAD_PJ_556_data_0) & "outputs: " & " LOAD_PJ_556_wire= "  & Convert_SLV_To_Hex_String(LOAD_PJ_556_wire));
      --
    end process; 
    -- equivalence LOAD_PJ_556_gather_scatter
    process(LOAD_PJ_556_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_PJ_556_data_0;
      ov(15 downto 0) := iv;
      LOAD_PJ_556_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator LOAD_ZJ_357_gather_scatter flow-through 
    process(LOAD_ZJ_357_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_ZJ_357_gather_scatter:flowthrough  inputs: " & " LOAD_ZJ_357_data_0 = "& Convert_SLV_To_Hex_String(LOAD_ZJ_357_data_0) & "outputs: " & " LOAD_ZJ_357_wire= "  & Convert_SLV_To_Hex_String(LOAD_ZJ_357_wire));
      --
    end process; 
    -- equivalence LOAD_ZJ_357_gather_scatter
    process(LOAD_ZJ_357_data_0) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(11 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_ZJ_357_data_0;
      ov(11 downto 0) := iv;
      LOAD_ZJ_357_wire <= ov(11 downto 0);
      --
    end process;
    -- logger for operator LOAD_one_366_gather_scatter flow-through 
    process(LOAD_one_366_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_one_366_gather_scatter:flowthrough  inputs: " & " LOAD_one_366_data_0 = "& Convert_SLV_To_Hex_String(LOAD_one_366_data_0) & "outputs: " & " LOAD_one_366_wire= "  & Convert_SLV_To_Hex_String(LOAD_one_366_wire));
      --
    end process; 
    -- equivalence LOAD_one_366_gather_scatter
    process(LOAD_one_366_data_0) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_one_366_data_0;
      ov(0 downto 0) := iv;
      LOAD_one_366_wire <= ov(0 downto 0);
      --
    end process;
    -- logger for operator LOAD_one_475_gather_scatter flow-through 
    process(LOAD_one_475_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_one_475_gather_scatter:flowthrough  inputs: " & " LOAD_one_475_data_0 = "& Convert_SLV_To_Hex_String(LOAD_one_475_data_0) & "outputs: " & " LOAD_one_475_wire= "  & Convert_SLV_To_Hex_String(LOAD_one_475_wire));
      --
    end process; 
    -- equivalence LOAD_one_475_gather_scatter
    process(LOAD_one_475_data_0) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_one_475_data_0;
      ov(0 downto 0) := iv;
      LOAD_one_475_wire <= ov(0 downto 0);
      --
    end process;
    -- logger for operator LOAD_total_603_gather_scatter flow-through 
    process(LOAD_total_603_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_total_603_gather_scatter:flowthrough  inputs: " & " LOAD_total_603_data_0 = "& Convert_SLV_To_Hex_String(LOAD_total_603_data_0) & "outputs: " & " LOAD_total_603_wire= "  & Convert_SLV_To_Hex_String(LOAD_total_603_wire));
      --
    end process; 
    -- equivalence LOAD_total_603_gather_scatter
    process(LOAD_total_603_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_total_603_data_0;
      ov(15 downto 0) := iv;
      LOAD_total_603_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator LOAD_total_622_gather_scatter flow-through 
    process(LOAD_total_622_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_total_622_gather_scatter:flowthrough  inputs: " & " LOAD_total_622_data_0 = "& Convert_SLV_To_Hex_String(LOAD_total_622_data_0) & "outputs: " & " LOAD_total_622_wire= "  & Convert_SLV_To_Hex_String(LOAD_total_622_wire));
      --
    end process; 
    -- equivalence LOAD_total_622_gather_scatter
    process(LOAD_total_622_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_total_622_data_0;
      ov(15 downto 0) := iv;
      LOAD_total_622_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator LOAD_zer_626_gather_scatter flow-through 
    process(LOAD_zer_626_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_zer_626_gather_scatter:flowthrough  inputs: " & " LOAD_zer_626_data_0 = "& Convert_SLV_To_Hex_String(LOAD_zer_626_data_0) & "outputs: " & " LOAD_zer_626_wire= "  & Convert_SLV_To_Hex_String(LOAD_zer_626_wire));
      --
    end process; 
    -- equivalence LOAD_zer_626_gather_scatter
    process(LOAD_zer_626_data_0) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_zer_626_data_0;
      ov(3 downto 0) := iv;
      LOAD_zer_626_wire <= ov(3 downto 0);
      --
    end process;
    -- logger for operator STORE_PJ_451_gather_scatter flow-through 
    process(STORE_PJ_451_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:STORE_PJ_451_gather_scatter:flowthrough  inputs: " & " konst_452_wire_constant = "& Convert_SLV_To_Hex_String(konst_452_wire_constant) & "outputs: " & " STORE_PJ_451_data_0= "  & Convert_SLV_To_Hex_String(STORE_PJ_451_data_0));
      --
    end process; 
    -- equivalence STORE_PJ_451_gather_scatter
    process(konst_452_wire_constant) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := konst_452_wire_constant;
      ov(15 downto 0) := iv;
      STORE_PJ_451_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator STORE_PJ_555_gather_scatter flow-through 
    process(STORE_PJ_555_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:STORE_PJ_555_gather_scatter:flowthrough  inputs: " & " ADD_u16_u16_558_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_558_wire) & "outputs: " & " STORE_PJ_555_data_0= "  & Convert_SLV_To_Hex_String(STORE_PJ_555_data_0));
      --
    end process; 
    -- equivalence STORE_PJ_555_gather_scatter
    process(ADD_u16_u16_558_wire) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u16_u16_558_wire;
      ov(15 downto 0) := iv;
      STORE_PJ_555_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator STORE_total_573_gather_scatter flow-through 
    process(STORE_total_573_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:STORE_total_573_gather_scatter:flowthrough  inputs: " & " konst_574_wire_constant = "& Convert_SLV_To_Hex_String(konst_574_wire_constant) & "outputs: " & " STORE_total_573_data_0= "  & Convert_SLV_To_Hex_String(STORE_total_573_data_0));
      --
    end process; 
    -- equivalence STORE_total_573_gather_scatter
    process(konst_574_wire_constant) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := konst_574_wire_constant;
      ov(15 downto 0) := iv;
      STORE_total_573_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator STORE_total_602_gather_scatter flow-through 
    process(STORE_total_602_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:STORE_total_602_gather_scatter:flowthrough  inputs: " & " ADD_u16_u16_606_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_606_wire) & "outputs: " & " STORE_total_602_data_0= "  & Convert_SLV_To_Hex_String(STORE_total_602_data_0));
      --
    end process; 
    -- equivalence STORE_total_602_gather_scatter
    process(ADD_u16_u16_606_wire) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u16_u16_606_wire;
      ov(15 downto 0) := iv;
      STORE_total_602_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_391_addr_0 flow-through 
    process(array_obj_ref_391_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_391_addr_0:flowthrough  inputs: " & " array_obj_ref_391_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_391_root_address) & "outputs: " & " array_obj_ref_391_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_391_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_391_addr_0
    process(array_obj_ref_391_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_391_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_391_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_391_gather_scatter flow-through 
    process(array_obj_ref_391_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_391_gather_scatter:flowthrough  inputs: " & " rdatak0_381 = "& Convert_SLV_To_Hex_String(rdatak0_381) & "outputs: " & " array_obj_ref_391_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_391_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_391_gather_scatter
    process(rdatak0_381) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdatak0_381;
      ov(15 downto 0) := iv;
      array_obj_ref_391_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_391_index_0_rename flow-through 
    process(R_T_341_delayed_12_0_390_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_391_index_0_rename:flowthrough  inputs: " & " R_T_341_delayed_12_0_390_resized = "& Convert_SLV_To_Hex_String(R_T_341_delayed_12_0_390_resized) & "outputs: " & " R_T_341_delayed_12_0_390_scaled= "  & Convert_SLV_To_Hex_String(R_T_341_delayed_12_0_390_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_391_index_0_rename
    process(R_T_341_delayed_12_0_390_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_T_341_delayed_12_0_390_resized;
      ov(3 downto 0) := iv;
      R_T_341_delayed_12_0_390_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_391_index_0_resize flow-through 
    process(R_T_341_delayed_12_0_390_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_391_index_0_resize:flowthrough  inputs: " & " T_341_delayed_12_0_389 = "& Convert_SLV_To_Hex_String(T_341_delayed_12_0_389) & "outputs: " & " R_T_341_delayed_12_0_390_resized= "  & Convert_SLV_To_Hex_String(R_T_341_delayed_12_0_390_resized));
      --
    end process; 
    -- equivalence array_obj_ref_391_index_0_resize
    process(T_341_delayed_12_0_389) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := T_341_delayed_12_0_389;
      ov := iv(3 downto 0);
      R_T_341_delayed_12_0_390_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_391_index_offset flow-through 
    process(array_obj_ref_391_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_391_index_offset:flowthrough  inputs: " & " R_T_341_delayed_12_0_390_scaled = "& Convert_SLV_To_Hex_String(R_T_341_delayed_12_0_390_scaled) & "outputs: " & " array_obj_ref_391_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_391_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_391_index_offset
    process(R_T_341_delayed_12_0_390_scaled) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_T_341_delayed_12_0_390_scaled;
      ov(3 downto 0) := iv;
      array_obj_ref_391_final_offset <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_391_root_address_inst flow-through 
    process(array_obj_ref_391_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_391_root_address_inst:flowthrough  inputs: " & " array_obj_ref_391_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_391_final_offset) & "outputs: " & " array_obj_ref_391_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_391_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_391_root_address_inst
    process(array_obj_ref_391_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_391_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_391_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_398_addr_0 flow-through 
    process(array_obj_ref_398_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_398_addr_0:flowthrough  inputs: " & " array_obj_ref_398_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_398_root_address) & "outputs: " & " array_obj_ref_398_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_398_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_398_addr_0
    process(array_obj_ref_398_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_398_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_398_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_398_gather_scatter flow-through 
    process(array_obj_ref_398_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_398_gather_scatter:flowthrough  inputs: " & " rdatak1_377 = "& Convert_SLV_To_Hex_String(rdatak1_377) & "outputs: " & " array_obj_ref_398_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_398_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_398_gather_scatter
    process(rdatak1_377) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdatak1_377;
      ov(15 downto 0) := iv;
      array_obj_ref_398_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_398_index_0_rename flow-through 
    process(R_TT_345_delayed_11_0_397_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_398_index_0_rename:flowthrough  inputs: " & " R_TT_345_delayed_11_0_397_resized = "& Convert_SLV_To_Hex_String(R_TT_345_delayed_11_0_397_resized) & "outputs: " & " R_TT_345_delayed_11_0_397_scaled= "  & Convert_SLV_To_Hex_String(R_TT_345_delayed_11_0_397_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_398_index_0_rename
    process(R_TT_345_delayed_11_0_397_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_TT_345_delayed_11_0_397_resized;
      ov(3 downto 0) := iv;
      R_TT_345_delayed_11_0_397_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_398_index_0_resize flow-through 
    process(R_TT_345_delayed_11_0_397_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_398_index_0_resize:flowthrough  inputs: " & " TT_345_delayed_11_0_396 = "& Convert_SLV_To_Hex_String(TT_345_delayed_11_0_396) & "outputs: " & " R_TT_345_delayed_11_0_397_resized= "  & Convert_SLV_To_Hex_String(R_TT_345_delayed_11_0_397_resized));
      --
    end process; 
    -- equivalence array_obj_ref_398_index_0_resize
    process(TT_345_delayed_11_0_396) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := TT_345_delayed_11_0_396;
      ov := iv(3 downto 0);
      R_TT_345_delayed_11_0_397_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_398_index_offset flow-through 
    process(array_obj_ref_398_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_398_index_offset:flowthrough  inputs: " & " R_TT_345_delayed_11_0_397_scaled = "& Convert_SLV_To_Hex_String(R_TT_345_delayed_11_0_397_scaled) & "outputs: " & " array_obj_ref_398_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_398_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_398_index_offset
    process(R_TT_345_delayed_11_0_397_scaled) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_TT_345_delayed_11_0_397_scaled;
      ov(3 downto 0) := iv;
      array_obj_ref_398_final_offset <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_398_root_address_inst flow-through 
    process(array_obj_ref_398_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_398_root_address_inst:flowthrough  inputs: " & " array_obj_ref_398_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_398_final_offset) & "outputs: " & " array_obj_ref_398_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_398_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_398_root_address_inst
    process(array_obj_ref_398_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_398_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_398_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_423_addr_0 flow-through 
    process(array_obj_ref_423_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_423_addr_0:flowthrough  inputs: " & " array_obj_ref_423_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_423_root_address) & "outputs: " & " array_obj_ref_423_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_423_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_423_addr_0
    process(array_obj_ref_423_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_423_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_423_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_423_gather_scatter flow-through 
    process(array_obj_ref_423_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_423_gather_scatter:flowthrough  inputs: " & " rdatak2_408 = "& Convert_SLV_To_Hex_String(rdatak2_408) & "outputs: " & " array_obj_ref_423_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_423_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_423_gather_scatter
    process(rdatak2_408) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdatak2_408;
      ov(15 downto 0) := iv;
      array_obj_ref_423_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_423_index_0_rename flow-through 
    process(R_TTT_367_delayed_11_0_422_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_423_index_0_rename:flowthrough  inputs: " & " R_TTT_367_delayed_11_0_422_resized = "& Convert_SLV_To_Hex_String(R_TTT_367_delayed_11_0_422_resized) & "outputs: " & " R_TTT_367_delayed_11_0_422_scaled= "  & Convert_SLV_To_Hex_String(R_TTT_367_delayed_11_0_422_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_423_index_0_rename
    process(R_TTT_367_delayed_11_0_422_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_TTT_367_delayed_11_0_422_resized;
      ov(3 downto 0) := iv;
      R_TTT_367_delayed_11_0_422_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_423_index_0_resize flow-through 
    process(R_TTT_367_delayed_11_0_422_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_423_index_0_resize:flowthrough  inputs: " & " TTT_367_delayed_11_0_421 = "& Convert_SLV_To_Hex_String(TTT_367_delayed_11_0_421) & "outputs: " & " R_TTT_367_delayed_11_0_422_resized= "  & Convert_SLV_To_Hex_String(R_TTT_367_delayed_11_0_422_resized));
      --
    end process; 
    -- equivalence array_obj_ref_423_index_0_resize
    process(TTT_367_delayed_11_0_421) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := TTT_367_delayed_11_0_421;
      ov := iv(3 downto 0);
      R_TTT_367_delayed_11_0_422_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_423_index_offset flow-through 
    process(array_obj_ref_423_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_423_index_offset:flowthrough  inputs: " & " R_TTT_367_delayed_11_0_422_scaled = "& Convert_SLV_To_Hex_String(R_TTT_367_delayed_11_0_422_scaled) & "outputs: " & " array_obj_ref_423_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_423_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_423_index_offset
    process(R_TTT_367_delayed_11_0_422_scaled) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_TTT_367_delayed_11_0_422_scaled;
      ov(3 downto 0) := iv;
      array_obj_ref_423_final_offset <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_423_root_address_inst flow-through 
    process(array_obj_ref_423_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_423_root_address_inst:flowthrough  inputs: " & " array_obj_ref_423_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_423_final_offset) & "outputs: " & " array_obj_ref_423_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_423_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_423_root_address_inst
    process(array_obj_ref_423_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_423_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_423_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_430_addr_0 flow-through 
    process(array_obj_ref_430_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_430_addr_0:flowthrough  inputs: " & " array_obj_ref_430_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_430_root_address) & "outputs: " & " array_obj_ref_430_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_430_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_430_addr_0
    process(array_obj_ref_430_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_430_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_430_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_430_gather_scatter flow-through 
    process(array_obj_ref_430_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_430_gather_scatter:flowthrough  inputs: " & " rdatak3_404 = "& Convert_SLV_To_Hex_String(rdatak3_404) & "outputs: " & " array_obj_ref_430_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_430_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_430_gather_scatter
    process(rdatak3_404) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdatak3_404;
      ov(15 downto 0) := iv;
      array_obj_ref_430_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_430_index_0_rename flow-through 
    process(R_TTTT_371_delayed_11_0_429_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_430_index_0_rename:flowthrough  inputs: " & " R_TTTT_371_delayed_11_0_429_resized = "& Convert_SLV_To_Hex_String(R_TTTT_371_delayed_11_0_429_resized) & "outputs: " & " R_TTTT_371_delayed_11_0_429_scaled= "  & Convert_SLV_To_Hex_String(R_TTTT_371_delayed_11_0_429_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_430_index_0_rename
    process(R_TTTT_371_delayed_11_0_429_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_TTTT_371_delayed_11_0_429_resized;
      ov(3 downto 0) := iv;
      R_TTTT_371_delayed_11_0_429_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_430_index_0_resize flow-through 
    process(R_TTTT_371_delayed_11_0_429_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_430_index_0_resize:flowthrough  inputs: " & " TTTT_371_delayed_11_0_428 = "& Convert_SLV_To_Hex_String(TTTT_371_delayed_11_0_428) & "outputs: " & " R_TTTT_371_delayed_11_0_429_resized= "  & Convert_SLV_To_Hex_String(R_TTTT_371_delayed_11_0_429_resized));
      --
    end process; 
    -- equivalence array_obj_ref_430_index_0_resize
    process(TTTT_371_delayed_11_0_428) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := TTTT_371_delayed_11_0_428;
      ov := iv(3 downto 0);
      R_TTTT_371_delayed_11_0_429_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_430_index_offset flow-through 
    process(array_obj_ref_430_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_430_index_offset:flowthrough  inputs: " & " R_TTTT_371_delayed_11_0_429_scaled = "& Convert_SLV_To_Hex_String(R_TTTT_371_delayed_11_0_429_scaled) & "outputs: " & " array_obj_ref_430_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_430_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_430_index_offset
    process(R_TTTT_371_delayed_11_0_429_scaled) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_TTTT_371_delayed_11_0_429_scaled;
      ov(3 downto 0) := iv;
      array_obj_ref_430_final_offset <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_430_root_address_inst flow-through 
    process(array_obj_ref_430_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_430_root_address_inst:flowthrough  inputs: " & " array_obj_ref_430_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_430_final_offset) & "outputs: " & " array_obj_ref_430_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_430_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_430_root_address_inst
    process(array_obj_ref_430_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_430_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_430_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_508_addr_0 flow-through 
    process(array_obj_ref_508_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_508_addr_0:flowthrough  inputs: " & " array_obj_ref_508_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_508_root_address) & "outputs: " & " array_obj_ref_508_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_508_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_508_addr_0
    process(array_obj_ref_508_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_508_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_508_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_508_gather_scatter flow-through 
    process(array_obj_ref_508_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_508_gather_scatter:flowthrough  inputs: " & " rdatai0_498 = "& Convert_SLV_To_Hex_String(rdatai0_498) & "outputs: " & " array_obj_ref_508_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_508_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_508_gather_scatter
    process(rdatai0_498) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdatai0_498;
      ov(15 downto 0) := iv;
      array_obj_ref_508_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_508_index_0_rename flow-through 
    process(R_PJ_440_delayed_7_0_507_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_508_index_0_rename:flowthrough  inputs: " & " R_PJ_440_delayed_7_0_507_resized = "& Convert_SLV_To_Hex_String(R_PJ_440_delayed_7_0_507_resized) & "outputs: " & " R_PJ_440_delayed_7_0_507_scaled= "  & Convert_SLV_To_Hex_String(R_PJ_440_delayed_7_0_507_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_508_index_0_rename
    process(R_PJ_440_delayed_7_0_507_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_PJ_440_delayed_7_0_507_resized;
      ov(3 downto 0) := iv;
      R_PJ_440_delayed_7_0_507_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_508_index_0_resize flow-through 
    process(R_PJ_440_delayed_7_0_507_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_508_index_0_resize:flowthrough  inputs: " & " PJ_440_delayed_7_0_506 = "& Convert_SLV_To_Hex_String(PJ_440_delayed_7_0_506) & "outputs: " & " R_PJ_440_delayed_7_0_507_resized= "  & Convert_SLV_To_Hex_String(R_PJ_440_delayed_7_0_507_resized));
      --
    end process; 
    -- equivalence array_obj_ref_508_index_0_resize
    process(PJ_440_delayed_7_0_506) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := PJ_440_delayed_7_0_506;
      ov := iv(3 downto 0);
      R_PJ_440_delayed_7_0_507_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_508_index_offset flow-through 
    process(array_obj_ref_508_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_508_index_offset:flowthrough  inputs: " & " R_PJ_440_delayed_7_0_507_scaled = "& Convert_SLV_To_Hex_String(R_PJ_440_delayed_7_0_507_scaled) & "outputs: " & " array_obj_ref_508_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_508_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_508_index_offset
    process(R_PJ_440_delayed_7_0_507_scaled) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_PJ_440_delayed_7_0_507_scaled;
      ov(3 downto 0) := iv;
      array_obj_ref_508_final_offset <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_508_root_address_inst flow-through 
    process(array_obj_ref_508_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_508_root_address_inst:flowthrough  inputs: " & " array_obj_ref_508_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_508_final_offset) & "outputs: " & " array_obj_ref_508_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_508_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_508_root_address_inst
    process(array_obj_ref_508_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_508_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_508_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_515_addr_0 flow-through 
    process(array_obj_ref_515_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_515_addr_0:flowthrough  inputs: " & " array_obj_ref_515_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_515_root_address) & "outputs: " & " array_obj_ref_515_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_515_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_515_addr_0
    process(array_obj_ref_515_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_515_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_515_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_515_gather_scatter flow-through 
    process(array_obj_ref_515_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_515_gather_scatter:flowthrough  inputs: " & " rdatai1_494 = "& Convert_SLV_To_Hex_String(rdatai1_494) & "outputs: " & " array_obj_ref_515_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_515_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_515_gather_scatter
    process(rdatai1_494) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdatai1_494;
      ov(15 downto 0) := iv;
      array_obj_ref_515_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_515_index_0_rename flow-through 
    process(R_PPJ_444_delayed_6_0_514_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_515_index_0_rename:flowthrough  inputs: " & " R_PPJ_444_delayed_6_0_514_resized = "& Convert_SLV_To_Hex_String(R_PPJ_444_delayed_6_0_514_resized) & "outputs: " & " R_PPJ_444_delayed_6_0_514_scaled= "  & Convert_SLV_To_Hex_String(R_PPJ_444_delayed_6_0_514_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_515_index_0_rename
    process(R_PPJ_444_delayed_6_0_514_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_PPJ_444_delayed_6_0_514_resized;
      ov(3 downto 0) := iv;
      R_PPJ_444_delayed_6_0_514_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_515_index_0_resize flow-through 
    process(R_PPJ_444_delayed_6_0_514_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_515_index_0_resize:flowthrough  inputs: " & " PPJ_444_delayed_6_0_513 = "& Convert_SLV_To_Hex_String(PPJ_444_delayed_6_0_513) & "outputs: " & " R_PPJ_444_delayed_6_0_514_resized= "  & Convert_SLV_To_Hex_String(R_PPJ_444_delayed_6_0_514_resized));
      --
    end process; 
    -- equivalence array_obj_ref_515_index_0_resize
    process(PPJ_444_delayed_6_0_513) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := PPJ_444_delayed_6_0_513;
      ov := iv(3 downto 0);
      R_PPJ_444_delayed_6_0_514_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_515_index_offset flow-through 
    process(array_obj_ref_515_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_515_index_offset:flowthrough  inputs: " & " R_PPJ_444_delayed_6_0_514_scaled = "& Convert_SLV_To_Hex_String(R_PPJ_444_delayed_6_0_514_scaled) & "outputs: " & " array_obj_ref_515_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_515_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_515_index_offset
    process(R_PPJ_444_delayed_6_0_514_scaled) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_PPJ_444_delayed_6_0_514_scaled;
      ov(3 downto 0) := iv;
      array_obj_ref_515_final_offset <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_515_root_address_inst flow-through 
    process(array_obj_ref_515_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_515_root_address_inst:flowthrough  inputs: " & " array_obj_ref_515_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_515_final_offset) & "outputs: " & " array_obj_ref_515_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_515_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_515_root_address_inst
    process(array_obj_ref_515_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_515_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_515_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_540_addr_0 flow-through 
    process(array_obj_ref_540_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_540_addr_0:flowthrough  inputs: " & " array_obj_ref_540_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_540_root_address) & "outputs: " & " array_obj_ref_540_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_540_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_540_addr_0
    process(array_obj_ref_540_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_540_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_540_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_540_gather_scatter flow-through 
    process(array_obj_ref_540_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_540_gather_scatter:flowthrough  inputs: " & " rdatai2_525 = "& Convert_SLV_To_Hex_String(rdatai2_525) & "outputs: " & " array_obj_ref_540_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_540_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_540_gather_scatter
    process(rdatai2_525) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdatai2_525;
      ov(15 downto 0) := iv;
      array_obj_ref_540_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_540_index_0_rename flow-through 
    process(R_PPPJ_466_delayed_6_0_539_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_540_index_0_rename:flowthrough  inputs: " & " R_PPPJ_466_delayed_6_0_539_resized = "& Convert_SLV_To_Hex_String(R_PPPJ_466_delayed_6_0_539_resized) & "outputs: " & " R_PPPJ_466_delayed_6_0_539_scaled= "  & Convert_SLV_To_Hex_String(R_PPPJ_466_delayed_6_0_539_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_540_index_0_rename
    process(R_PPPJ_466_delayed_6_0_539_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_PPPJ_466_delayed_6_0_539_resized;
      ov(3 downto 0) := iv;
      R_PPPJ_466_delayed_6_0_539_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_540_index_0_resize flow-through 
    process(R_PPPJ_466_delayed_6_0_539_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_540_index_0_resize:flowthrough  inputs: " & " PPPJ_466_delayed_6_0_538 = "& Convert_SLV_To_Hex_String(PPPJ_466_delayed_6_0_538) & "outputs: " & " R_PPPJ_466_delayed_6_0_539_resized= "  & Convert_SLV_To_Hex_String(R_PPPJ_466_delayed_6_0_539_resized));
      --
    end process; 
    -- equivalence array_obj_ref_540_index_0_resize
    process(PPPJ_466_delayed_6_0_538) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := PPPJ_466_delayed_6_0_538;
      ov := iv(3 downto 0);
      R_PPPJ_466_delayed_6_0_539_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_540_index_offset flow-through 
    process(array_obj_ref_540_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_540_index_offset:flowthrough  inputs: " & " R_PPPJ_466_delayed_6_0_539_scaled = "& Convert_SLV_To_Hex_String(R_PPPJ_466_delayed_6_0_539_scaled) & "outputs: " & " array_obj_ref_540_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_540_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_540_index_offset
    process(R_PPPJ_466_delayed_6_0_539_scaled) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_PPPJ_466_delayed_6_0_539_scaled;
      ov(3 downto 0) := iv;
      array_obj_ref_540_final_offset <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_540_root_address_inst flow-through 
    process(array_obj_ref_540_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_540_root_address_inst:flowthrough  inputs: " & " array_obj_ref_540_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_540_final_offset) & "outputs: " & " array_obj_ref_540_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_540_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_540_root_address_inst
    process(array_obj_ref_540_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_540_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_540_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_547_addr_0 flow-through 
    process(array_obj_ref_547_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_547_addr_0:flowthrough  inputs: " & " array_obj_ref_547_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_547_root_address) & "outputs: " & " array_obj_ref_547_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_547_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_547_addr_0
    process(array_obj_ref_547_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_547_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_547_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_547_gather_scatter flow-through 
    process(array_obj_ref_547_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_547_gather_scatter:flowthrough  inputs: " & " rdatai3_521 = "& Convert_SLV_To_Hex_String(rdatai3_521) & "outputs: " & " array_obj_ref_547_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_547_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_547_gather_scatter
    process(rdatai3_521) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdatai3_521;
      ov(15 downto 0) := iv;
      array_obj_ref_547_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_547_index_0_rename flow-through 
    process(R_PPPPJ_470_delayed_6_0_546_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_547_index_0_rename:flowthrough  inputs: " & " R_PPPPJ_470_delayed_6_0_546_resized = "& Convert_SLV_To_Hex_String(R_PPPPJ_470_delayed_6_0_546_resized) & "outputs: " & " R_PPPPJ_470_delayed_6_0_546_scaled= "  & Convert_SLV_To_Hex_String(R_PPPPJ_470_delayed_6_0_546_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_547_index_0_rename
    process(R_PPPPJ_470_delayed_6_0_546_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_PPPPJ_470_delayed_6_0_546_resized;
      ov(3 downto 0) := iv;
      R_PPPPJ_470_delayed_6_0_546_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_547_index_0_resize flow-through 
    process(R_PPPPJ_470_delayed_6_0_546_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_547_index_0_resize:flowthrough  inputs: " & " PPPPJ_470_delayed_6_0_545 = "& Convert_SLV_To_Hex_String(PPPPJ_470_delayed_6_0_545) & "outputs: " & " R_PPPPJ_470_delayed_6_0_546_resized= "  & Convert_SLV_To_Hex_String(R_PPPPJ_470_delayed_6_0_546_resized));
      --
    end process; 
    -- equivalence array_obj_ref_547_index_0_resize
    process(PPPPJ_470_delayed_6_0_545) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := PPPPJ_470_delayed_6_0_545;
      ov := iv(3 downto 0);
      R_PPPPJ_470_delayed_6_0_546_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_547_index_offset flow-through 
    process(array_obj_ref_547_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_547_index_offset:flowthrough  inputs: " & " R_PPPPJ_470_delayed_6_0_546_scaled = "& Convert_SLV_To_Hex_String(R_PPPPJ_470_delayed_6_0_546_scaled) & "outputs: " & " array_obj_ref_547_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_547_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_547_index_offset
    process(R_PPPPJ_470_delayed_6_0_546_scaled) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_PPPPJ_470_delayed_6_0_546_scaled;
      ov(3 downto 0) := iv;
      array_obj_ref_547_final_offset <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_547_root_address_inst flow-through 
    process(array_obj_ref_547_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_547_root_address_inst:flowthrough  inputs: " & " array_obj_ref_547_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_547_final_offset) & "outputs: " & " array_obj_ref_547_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_547_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_547_root_address_inst
    process(array_obj_ref_547_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_547_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_547_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_587_addr_0 flow-through 
    process(array_obj_ref_587_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_587_addr_0:flowthrough  inputs: " & " array_obj_ref_587_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_587_root_address) & "outputs: " & " array_obj_ref_587_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_587_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_587_addr_0
    process(array_obj_ref_587_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_587_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_587_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_587_gather_scatter flow-through 
    process(imag1_588) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_587_gather_scatter:flowthrough  inputs: " & " array_obj_ref_587_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_587_data_0) & "outputs: " & " imag1_588= "  & Convert_SLV_To_Hex_String(imag1_588));
      --
    end process; 
    -- equivalence array_obj_ref_587_gather_scatter
    process(array_obj_ref_587_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_587_data_0;
      ov(15 downto 0) := iv;
      imag1_588 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_587_index_0_rename flow-through 
    process(R_K_586_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_587_index_0_rename:flowthrough  inputs: " & " R_K_586_resized = "& Convert_SLV_To_Hex_String(R_K_586_resized) & "outputs: " & " R_K_586_scaled= "  & Convert_SLV_To_Hex_String(R_K_586_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_587_index_0_rename
    process(R_K_586_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_K_586_resized;
      ov(3 downto 0) := iv;
      R_K_586_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_587_index_0_resize flow-through 
    process(R_K_586_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_587_index_0_resize:flowthrough  inputs: " & " K_579 = "& Convert_SLV_To_Hex_String(K_579) & "outputs: " & " R_K_586_resized= "  & Convert_SLV_To_Hex_String(R_K_586_resized));
      --
    end process; 
    -- equivalence array_obj_ref_587_index_0_resize
    process(K_579) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := K_579;
      ov := iv(3 downto 0);
      R_K_586_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_587_index_offset flow-through 
    process(array_obj_ref_587_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_587_index_offset:flowthrough  inputs: " & " R_K_586_scaled = "& Convert_SLV_To_Hex_String(R_K_586_scaled) & "outputs: " & " array_obj_ref_587_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_587_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_587_index_offset
    process(R_K_586_scaled) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_K_586_scaled;
      ov(3 downto 0) := iv;
      array_obj_ref_587_final_offset <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_587_root_address_inst flow-through 
    process(array_obj_ref_587_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_587_root_address_inst:flowthrough  inputs: " & " array_obj_ref_587_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_587_final_offset) & "outputs: " & " array_obj_ref_587_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_587_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_587_root_address_inst
    process(array_obj_ref_587_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_587_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_587_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_591_addr_0 flow-through 
    process(array_obj_ref_591_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_591_addr_0:flowthrough  inputs: " & " array_obj_ref_591_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_591_root_address) & "outputs: " & " array_obj_ref_591_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_591_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_591_addr_0
    process(array_obj_ref_591_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_591_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_591_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_591_gather_scatter flow-through 
    process(ker1_592) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_591_gather_scatter:flowthrough  inputs: " & " array_obj_ref_591_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_591_data_0) & "outputs: " & " ker1_592= "  & Convert_SLV_To_Hex_String(ker1_592));
      --
    end process; 
    -- equivalence array_obj_ref_591_gather_scatter
    process(array_obj_ref_591_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_591_data_0;
      ov(15 downto 0) := iv;
      ker1_592 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_591_index_0_rename flow-through 
    process(R_K_590_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_591_index_0_rename:flowthrough  inputs: " & " R_K_590_resized = "& Convert_SLV_To_Hex_String(R_K_590_resized) & "outputs: " & " R_K_590_scaled= "  & Convert_SLV_To_Hex_String(R_K_590_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_591_index_0_rename
    process(R_K_590_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_K_590_resized;
      ov(3 downto 0) := iv;
      R_K_590_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_591_index_0_resize flow-through 
    process(R_K_590_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_591_index_0_resize:flowthrough  inputs: " & " K_579 = "& Convert_SLV_To_Hex_String(K_579) & "outputs: " & " R_K_590_resized= "  & Convert_SLV_To_Hex_String(R_K_590_resized));
      --
    end process; 
    -- equivalence array_obj_ref_591_index_0_resize
    process(K_579) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := K_579;
      ov := iv(3 downto 0);
      R_K_590_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_591_index_offset flow-through 
    process(array_obj_ref_591_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_591_index_offset:flowthrough  inputs: " & " R_K_590_scaled = "& Convert_SLV_To_Hex_String(R_K_590_scaled) & "outputs: " & " array_obj_ref_591_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_591_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_591_index_offset
    process(R_K_590_scaled) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_K_590_scaled;
      ov(3 downto 0) := iv;
      array_obj_ref_591_final_offset <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_591_root_address_inst flow-through 
    process(array_obj_ref_591_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_591_root_address_inst:flowthrough  inputs: " & " array_obj_ref_591_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_591_final_offset) & "outputs: " & " array_obj_ref_591_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_591_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_591_root_address_inst
    process(array_obj_ref_591_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_591_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_591_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_597_addr_0 flow-through 
    process(array_obj_ref_597_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_597_addr_0:flowthrough  inputs: " & " array_obj_ref_597_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_597_root_address) & "outputs: " & " array_obj_ref_597_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_597_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_597_addr_0
    process(array_obj_ref_597_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_597_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_597_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_597_gather_scatter flow-through 
    process(array_obj_ref_597_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_597_gather_scatter:flowthrough  inputs: " & " MUL_u16_u16_600_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_600_wire) & "outputs: " & " array_obj_ref_597_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_597_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_597_gather_scatter
    process(MUL_u16_u16_600_wire) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := MUL_u16_u16_600_wire;
      ov(15 downto 0) := iv;
      array_obj_ref_597_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_597_index_0_rename flow-through 
    process(R_K_517_delayed_5_0_596_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_597_index_0_rename:flowthrough  inputs: " & " R_K_517_delayed_5_0_596_resized = "& Convert_SLV_To_Hex_String(R_K_517_delayed_5_0_596_resized) & "outputs: " & " R_K_517_delayed_5_0_596_scaled= "  & Convert_SLV_To_Hex_String(R_K_517_delayed_5_0_596_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_597_index_0_rename
    process(R_K_517_delayed_5_0_596_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_K_517_delayed_5_0_596_resized;
      ov(3 downto 0) := iv;
      R_K_517_delayed_5_0_596_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_597_index_0_resize flow-through 
    process(R_K_517_delayed_5_0_596_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_597_index_0_resize:flowthrough  inputs: " & " K_517_delayed_5_0_595 = "& Convert_SLV_To_Hex_String(K_517_delayed_5_0_595) & "outputs: " & " R_K_517_delayed_5_0_596_resized= "  & Convert_SLV_To_Hex_String(R_K_517_delayed_5_0_596_resized));
      --
    end process; 
    -- equivalence array_obj_ref_597_index_0_resize
    process(K_517_delayed_5_0_595) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := K_517_delayed_5_0_595;
      ov := iv(3 downto 0);
      R_K_517_delayed_5_0_596_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_597_index_offset flow-through 
    process(array_obj_ref_597_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_597_index_offset:flowthrough  inputs: " & " R_K_517_delayed_5_0_596_scaled = "& Convert_SLV_To_Hex_String(R_K_517_delayed_5_0_596_scaled) & "outputs: " & " array_obj_ref_597_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_597_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_597_index_offset
    process(R_K_517_delayed_5_0_596_scaled) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_K_517_delayed_5_0_596_scaled;
      ov(3 downto 0) := iv;
      array_obj_ref_597_final_offset <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_597_root_address_inst flow-through 
    process(array_obj_ref_597_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_597_root_address_inst:flowthrough  inputs: " & " array_obj_ref_597_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_597_final_offset) & "outputs: " & " array_obj_ref_597_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_597_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_597_root_address_inst
    process(array_obj_ref_597_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_597_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_597_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_605_addr_0 flow-through 
    process(array_obj_ref_605_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_605_addr_0:flowthrough  inputs: " & " array_obj_ref_605_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_605_root_address) & "outputs: " & " array_obj_ref_605_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_605_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_605_addr_0
    process(array_obj_ref_605_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_605_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_605_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_605_gather_scatter flow-through 
    process(array_obj_ref_605_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_605_gather_scatter:flowthrough  inputs: " & " array_obj_ref_605_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_605_data_0) & "outputs: " & " array_obj_ref_605_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_605_wire));
      --
    end process; 
    -- equivalence array_obj_ref_605_gather_scatter
    process(array_obj_ref_605_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_605_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_605_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_605_index_0_rename flow-through 
    process(R_K_604_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_605_index_0_rename:flowthrough  inputs: " & " R_K_604_resized = "& Convert_SLV_To_Hex_String(R_K_604_resized) & "outputs: " & " R_K_604_scaled= "  & Convert_SLV_To_Hex_String(R_K_604_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_605_index_0_rename
    process(R_K_604_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_K_604_resized;
      ov(3 downto 0) := iv;
      R_K_604_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_605_index_0_resize flow-through 
    process(R_K_604_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_605_index_0_resize:flowthrough  inputs: " & " K_579 = "& Convert_SLV_To_Hex_String(K_579) & "outputs: " & " R_K_604_resized= "  & Convert_SLV_To_Hex_String(R_K_604_resized));
      --
    end process; 
    -- equivalence array_obj_ref_605_index_0_resize
    process(K_579) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := K_579;
      ov := iv(3 downto 0);
      R_K_604_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_605_index_offset flow-through 
    process(array_obj_ref_605_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_605_index_offset:flowthrough  inputs: " & " R_K_604_scaled = "& Convert_SLV_To_Hex_String(R_K_604_scaled) & "outputs: " & " array_obj_ref_605_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_605_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_605_index_offset
    process(R_K_604_scaled) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_K_604_scaled;
      ov(3 downto 0) := iv;
      array_obj_ref_605_final_offset <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_605_root_address_inst flow-through 
    process(array_obj_ref_605_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_605_root_address_inst:flowthrough  inputs: " & " array_obj_ref_605_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_605_final_offset) & "outputs: " & " array_obj_ref_605_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_605_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_605_root_address_inst
    process(array_obj_ref_605_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_605_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_605_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_637_addr_0 flow-through 
    process(array_obj_ref_637_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_637_addr_0:flowthrough  inputs: " & " array_obj_ref_637_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_637_root_address) & "outputs: " & " array_obj_ref_637_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_637_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_637_addr_0
    process(array_obj_ref_637_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_637_root_address;
      ov(10 downto 0) := iv;
      array_obj_ref_637_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_637_gather_scatter flow-through 
    process(array_obj_ref_637_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_637_gather_scatter:flowthrough  inputs: " & " array_obj_ref_637_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_637_data_0) & "outputs: " & " array_obj_ref_637_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_637_wire));
      --
    end process; 
    -- equivalence array_obj_ref_637_gather_scatter
    process(array_obj_ref_637_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_637_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_637_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_637_index_0_rename flow-through 
    process(R_f_636_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_637_index_0_rename:flowthrough  inputs: " & " R_f_636_resized = "& Convert_SLV_To_Hex_String(R_f_636_resized) & "outputs: " & " R_f_636_scaled= "  & Convert_SLV_To_Hex_String(R_f_636_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_637_index_0_rename
    process(R_f_636_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_f_636_resized;
      ov(10 downto 0) := iv;
      R_f_636_scaled <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_637_index_0_resize flow-through 
    process(R_f_636_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_637_index_0_resize:flowthrough  inputs: " & " f_631 = "& Convert_SLV_To_Hex_String(f_631) & "outputs: " & " R_f_636_resized= "  & Convert_SLV_To_Hex_String(R_f_636_resized));
      --
    end process; 
    -- equivalence array_obj_ref_637_index_0_resize
    process(f_631) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := f_631;
      ov := iv(10 downto 0);
      R_f_636_resized <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_637_index_offset flow-through 
    process(array_obj_ref_637_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_637_index_offset:flowthrough  inputs: " & " R_f_636_scaled = "& Convert_SLV_To_Hex_String(R_f_636_scaled) & "outputs: " & " array_obj_ref_637_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_637_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_637_index_offset
    process(R_f_636_scaled) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_f_636_scaled;
      ov(10 downto 0) := iv;
      array_obj_ref_637_final_offset <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_637_root_address_inst flow-through 
    process(array_obj_ref_637_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_637_root_address_inst:flowthrough  inputs: " & " array_obj_ref_637_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_637_final_offset) & "outputs: " & " array_obj_ref_637_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_637_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_637_root_address_inst
    process(array_obj_ref_637_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_637_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_637_root_address <= ov(10 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_657_addr_0 flow-through 
    process(array_obj_ref_657_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_657_addr_0:flowthrough  inputs: " & " array_obj_ref_657_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_657_root_address) & "outputs: " & " array_obj_ref_657_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_657_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_657_addr_0
    process(array_obj_ref_657_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_657_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_657_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_657_gather_scatter flow-through 
    process(array_obj_ref_657_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_657_gather_scatter:flowthrough  inputs: " & " array_obj_ref_659_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_659_wire) & "outputs: " & " array_obj_ref_657_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_657_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_657_gather_scatter
    process(array_obj_ref_659_wire) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_659_wire;
      ov(15 downto 0) := iv;
      array_obj_ref_657_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_657_index_0_rename flow-through 
    process(R_H_574_delayed_5_0_656_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_657_index_0_rename:flowthrough  inputs: " & " R_H_574_delayed_5_0_656_resized = "& Convert_SLV_To_Hex_String(R_H_574_delayed_5_0_656_resized) & "outputs: " & " R_H_574_delayed_5_0_656_scaled= "  & Convert_SLV_To_Hex_String(R_H_574_delayed_5_0_656_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_657_index_0_rename
    process(R_H_574_delayed_5_0_656_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_H_574_delayed_5_0_656_resized;
      ov(3 downto 0) := iv;
      R_H_574_delayed_5_0_656_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_657_index_0_resize flow-through 
    process(R_H_574_delayed_5_0_656_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_657_index_0_resize:flowthrough  inputs: " & " H_574_delayed_5_0_655 = "& Convert_SLV_To_Hex_String(H_574_delayed_5_0_655) & "outputs: " & " R_H_574_delayed_5_0_656_resized= "  & Convert_SLV_To_Hex_String(R_H_574_delayed_5_0_656_resized));
      --
    end process; 
    -- equivalence array_obj_ref_657_index_0_resize
    process(H_574_delayed_5_0_655) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := H_574_delayed_5_0_655;
      ov := iv(3 downto 0);
      R_H_574_delayed_5_0_656_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_657_index_offset flow-through 
    process(array_obj_ref_657_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_657_index_offset:flowthrough  inputs: " & " R_H_574_delayed_5_0_656_scaled = "& Convert_SLV_To_Hex_String(R_H_574_delayed_5_0_656_scaled) & "outputs: " & " array_obj_ref_657_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_657_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_657_index_offset
    process(R_H_574_delayed_5_0_656_scaled) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_H_574_delayed_5_0_656_scaled;
      ov(3 downto 0) := iv;
      array_obj_ref_657_final_offset <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_657_root_address_inst flow-through 
    process(array_obj_ref_657_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_657_root_address_inst:flowthrough  inputs: " & " array_obj_ref_657_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_657_final_offset) & "outputs: " & " array_obj_ref_657_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_657_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_657_root_address_inst
    process(array_obj_ref_657_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_657_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_657_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_659_addr_0 flow-through 
    process(array_obj_ref_659_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_659_addr_0:flowthrough  inputs: " & " array_obj_ref_659_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_659_root_address) & "outputs: " & " array_obj_ref_659_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_659_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_659_addr_0
    process(array_obj_ref_659_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_659_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_659_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_659_gather_scatter flow-through 
    process(array_obj_ref_659_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_659_gather_scatter:flowthrough  inputs: " & " array_obj_ref_659_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_659_data_0) & "outputs: " & " array_obj_ref_659_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_659_wire));
      --
    end process; 
    -- equivalence array_obj_ref_659_gather_scatter
    process(array_obj_ref_659_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_659_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_659_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_659_index_0_rename flow-through 
    process(R_HH_658_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_659_index_0_rename:flowthrough  inputs: " & " R_HH_658_resized = "& Convert_SLV_To_Hex_String(R_HH_658_resized) & "outputs: " & " R_HH_658_scaled= "  & Convert_SLV_To_Hex_String(R_HH_658_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_659_index_0_rename
    process(R_HH_658_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_HH_658_resized;
      ov(3 downto 0) := iv;
      R_HH_658_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_659_index_0_resize flow-through 
    process(R_HH_658_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_659_index_0_resize:flowthrough  inputs: " & " HH_652 = "& Convert_SLV_To_Hex_String(HH_652) & "outputs: " & " R_HH_658_resized= "  & Convert_SLV_To_Hex_String(R_HH_658_resized));
      --
    end process; 
    -- equivalence array_obj_ref_659_index_0_resize
    process(HH_652) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := HH_652;
      ov := iv(3 downto 0);
      R_HH_658_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_659_index_offset flow-through 
    process(array_obj_ref_659_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_659_index_offset:flowthrough  inputs: " & " R_HH_658_scaled = "& Convert_SLV_To_Hex_String(R_HH_658_scaled) & "outputs: " & " array_obj_ref_659_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_659_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_659_index_offset
    process(R_HH_658_scaled) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_HH_658_scaled;
      ov(3 downto 0) := iv;
      array_obj_ref_659_final_offset <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_659_root_address_inst flow-through 
    process(array_obj_ref_659_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_659_root_address_inst:flowthrough  inputs: " & " array_obj_ref_659_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_659_final_offset) & "outputs: " & " array_obj_ref_659_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_659_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_659_root_address_inst
    process(array_obj_ref_659_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_659_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_659_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_670_addr_0 flow-through 
    process(array_obj_ref_670_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_670_addr_0:flowthrough  inputs: " & " array_obj_ref_670_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_670_root_address) & "outputs: " & " array_obj_ref_670_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_670_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_670_addr_0
    process(array_obj_ref_670_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_670_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_670_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_670_gather_scatter flow-through 
    process(array_obj_ref_670_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_670_gather_scatter:flowthrough  inputs: " & " array_obj_ref_672_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_672_wire) & "outputs: " & " array_obj_ref_670_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_670_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_670_gather_scatter
    process(array_obj_ref_672_wire) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_672_wire;
      ov(15 downto 0) := iv;
      array_obj_ref_670_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_670_index_0_rename flow-through 
    process(R_HH_584_delayed_4_0_669_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_670_index_0_rename:flowthrough  inputs: " & " R_HH_584_delayed_4_0_669_resized = "& Convert_SLV_To_Hex_String(R_HH_584_delayed_4_0_669_resized) & "outputs: " & " R_HH_584_delayed_4_0_669_scaled= "  & Convert_SLV_To_Hex_String(R_HH_584_delayed_4_0_669_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_670_index_0_rename
    process(R_HH_584_delayed_4_0_669_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_HH_584_delayed_4_0_669_resized;
      ov(3 downto 0) := iv;
      R_HH_584_delayed_4_0_669_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_670_index_0_resize flow-through 
    process(R_HH_584_delayed_4_0_669_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_670_index_0_resize:flowthrough  inputs: " & " HH_584_delayed_4_0_668 = "& Convert_SLV_To_Hex_String(HH_584_delayed_4_0_668) & "outputs: " & " R_HH_584_delayed_4_0_669_resized= "  & Convert_SLV_To_Hex_String(R_HH_584_delayed_4_0_669_resized));
      --
    end process; 
    -- equivalence array_obj_ref_670_index_0_resize
    process(HH_584_delayed_4_0_668) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := HH_584_delayed_4_0_668;
      ov := iv(3 downto 0);
      R_HH_584_delayed_4_0_669_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_670_index_offset flow-through 
    process(array_obj_ref_670_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_670_index_offset:flowthrough  inputs: " & " R_HH_584_delayed_4_0_669_scaled = "& Convert_SLV_To_Hex_String(R_HH_584_delayed_4_0_669_scaled) & "outputs: " & " array_obj_ref_670_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_670_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_670_index_offset
    process(R_HH_584_delayed_4_0_669_scaled) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_HH_584_delayed_4_0_669_scaled;
      ov(3 downto 0) := iv;
      array_obj_ref_670_final_offset <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_670_root_address_inst flow-through 
    process(array_obj_ref_670_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_670_root_address_inst:flowthrough  inputs: " & " array_obj_ref_670_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_670_final_offset) & "outputs: " & " array_obj_ref_670_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_670_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_670_root_address_inst
    process(array_obj_ref_670_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_670_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_670_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_672_addr_0 flow-through 
    process(array_obj_ref_672_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_672_addr_0:flowthrough  inputs: " & " array_obj_ref_672_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_672_root_address) & "outputs: " & " array_obj_ref_672_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_672_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_672_addr_0
    process(array_obj_ref_672_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_672_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_672_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_672_gather_scatter flow-through 
    process(array_obj_ref_672_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_672_gather_scatter:flowthrough  inputs: " & " array_obj_ref_672_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_672_data_0) & "outputs: " & " array_obj_ref_672_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_672_wire));
      --
    end process; 
    -- equivalence array_obj_ref_672_gather_scatter
    process(array_obj_ref_672_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_672_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_672_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_672_index_0_rename flow-through 
    process(R_HHH_671_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_672_index_0_rename:flowthrough  inputs: " & " R_HHH_671_resized = "& Convert_SLV_To_Hex_String(R_HHH_671_resized) & "outputs: " & " R_HHH_671_scaled= "  & Convert_SLV_To_Hex_String(R_HHH_671_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_672_index_0_rename
    process(R_HHH_671_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_HHH_671_resized;
      ov(3 downto 0) := iv;
      R_HHH_671_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_672_index_0_resize flow-through 
    process(R_HHH_671_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_672_index_0_resize:flowthrough  inputs: " & " HHH_665 = "& Convert_SLV_To_Hex_String(HHH_665) & "outputs: " & " R_HHH_671_resized= "  & Convert_SLV_To_Hex_String(R_HHH_671_resized));
      --
    end process; 
    -- equivalence array_obj_ref_672_index_0_resize
    process(HHH_665) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := HHH_665;
      ov := iv(3 downto 0);
      R_HHH_671_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_672_index_offset flow-through 
    process(array_obj_ref_672_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_672_index_offset:flowthrough  inputs: " & " R_HHH_671_scaled = "& Convert_SLV_To_Hex_String(R_HHH_671_scaled) & "outputs: " & " array_obj_ref_672_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_672_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_672_index_offset
    process(R_HHH_671_scaled) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_HHH_671_scaled;
      ov(3 downto 0) := iv;
      array_obj_ref_672_final_offset <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_672_root_address_inst flow-through 
    process(array_obj_ref_672_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_672_root_address_inst:flowthrough  inputs: " & " array_obj_ref_672_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_672_final_offset) & "outputs: " & " array_obj_ref_672_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_672_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_672_root_address_inst
    process(array_obj_ref_672_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_672_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_672_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_683_addr_0 flow-through 
    process(array_obj_ref_683_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_683_addr_0:flowthrough  inputs: " & " array_obj_ref_683_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_683_root_address) & "outputs: " & " array_obj_ref_683_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_683_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_683_addr_0
    process(array_obj_ref_683_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_683_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_683_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_683_gather_scatter flow-through 
    process(array_obj_ref_683_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_683_gather_scatter:flowthrough  inputs: " & " array_obj_ref_685_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_685_wire) & "outputs: " & " array_obj_ref_683_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_683_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_683_gather_scatter
    process(array_obj_ref_685_wire) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_685_wire;
      ov(15 downto 0) := iv;
      array_obj_ref_683_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_683_index_0_rename flow-through 
    process(R_HHH_594_delayed_4_0_682_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_683_index_0_rename:flowthrough  inputs: " & " R_HHH_594_delayed_4_0_682_resized = "& Convert_SLV_To_Hex_String(R_HHH_594_delayed_4_0_682_resized) & "outputs: " & " R_HHH_594_delayed_4_0_682_scaled= "  & Convert_SLV_To_Hex_String(R_HHH_594_delayed_4_0_682_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_683_index_0_rename
    process(R_HHH_594_delayed_4_0_682_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_HHH_594_delayed_4_0_682_resized;
      ov(3 downto 0) := iv;
      R_HHH_594_delayed_4_0_682_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_683_index_0_resize flow-through 
    process(R_HHH_594_delayed_4_0_682_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_683_index_0_resize:flowthrough  inputs: " & " HHH_594_delayed_4_0_681 = "& Convert_SLV_To_Hex_String(HHH_594_delayed_4_0_681) & "outputs: " & " R_HHH_594_delayed_4_0_682_resized= "  & Convert_SLV_To_Hex_String(R_HHH_594_delayed_4_0_682_resized));
      --
    end process; 
    -- equivalence array_obj_ref_683_index_0_resize
    process(HHH_594_delayed_4_0_681) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := HHH_594_delayed_4_0_681;
      ov := iv(3 downto 0);
      R_HHH_594_delayed_4_0_682_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_683_index_offset flow-through 
    process(array_obj_ref_683_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_683_index_offset:flowthrough  inputs: " & " R_HHH_594_delayed_4_0_682_scaled = "& Convert_SLV_To_Hex_String(R_HHH_594_delayed_4_0_682_scaled) & "outputs: " & " array_obj_ref_683_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_683_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_683_index_offset
    process(R_HHH_594_delayed_4_0_682_scaled) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_HHH_594_delayed_4_0_682_scaled;
      ov(3 downto 0) := iv;
      array_obj_ref_683_final_offset <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_683_root_address_inst flow-through 
    process(array_obj_ref_683_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_683_root_address_inst:flowthrough  inputs: " & " array_obj_ref_683_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_683_final_offset) & "outputs: " & " array_obj_ref_683_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_683_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_683_root_address_inst
    process(array_obj_ref_683_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_683_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_683_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_685_addr_0 flow-through 
    process(array_obj_ref_685_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_685_addr_0:flowthrough  inputs: " & " array_obj_ref_685_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_685_root_address) & "outputs: " & " array_obj_ref_685_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_685_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_685_addr_0
    process(array_obj_ref_685_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_685_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_685_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_685_gather_scatter flow-through 
    process(array_obj_ref_685_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_685_gather_scatter:flowthrough  inputs: " & " array_obj_ref_685_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_685_data_0) & "outputs: " & " array_obj_ref_685_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_685_wire));
      --
    end process; 
    -- equivalence array_obj_ref_685_gather_scatter
    process(array_obj_ref_685_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_685_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_685_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_685_index_0_rename flow-through 
    process(R_HHHH_684_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_685_index_0_rename:flowthrough  inputs: " & " R_HHHH_684_resized = "& Convert_SLV_To_Hex_String(R_HHHH_684_resized) & "outputs: " & " R_HHHH_684_scaled= "  & Convert_SLV_To_Hex_String(R_HHHH_684_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_685_index_0_rename
    process(R_HHHH_684_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_HHHH_684_resized;
      ov(3 downto 0) := iv;
      R_HHHH_684_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_685_index_0_resize flow-through 
    process(R_HHHH_684_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_685_index_0_resize:flowthrough  inputs: " & " HHHH_678 = "& Convert_SLV_To_Hex_String(HHHH_678) & "outputs: " & " R_HHHH_684_resized= "  & Convert_SLV_To_Hex_String(R_HHHH_684_resized));
      --
    end process; 
    -- equivalence array_obj_ref_685_index_0_resize
    process(HHHH_678) --
      variable iv : std_logic_vector(11 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := HHHH_678;
      ov := iv(3 downto 0);
      R_HHHH_684_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_685_index_offset flow-through 
    process(array_obj_ref_685_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_685_index_offset:flowthrough  inputs: " & " R_HHHH_684_scaled = "& Convert_SLV_To_Hex_String(R_HHHH_684_scaled) & "outputs: " & " array_obj_ref_685_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_685_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_685_index_offset
    process(R_HHHH_684_scaled) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_HHHH_684_scaled;
      ov(3 downto 0) := iv;
      array_obj_ref_685_final_offset <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_685_root_address_inst flow-through 
    process(array_obj_ref_685_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_685_root_address_inst:flowthrough  inputs: " & " array_obj_ref_685_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_685_final_offset) & "outputs: " & " array_obj_ref_685_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_685_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_685_root_address_inst
    process(array_obj_ref_685_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_685_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_685_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_707_gather_scatter flow-through 
    process(array_obj_ref_707_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_707_gather_scatter:flowthrough  inputs: " & " slice_709_wire = "& Convert_SLV_To_Hex_String(slice_709_wire) & "outputs: " & " array_obj_ref_707_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_707_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_707_gather_scatter
    process(slice_709_wire) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := slice_709_wire;
      ov(15 downto 0) := iv;
      array_obj_ref_707_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_712_gather_scatter flow-through 
    process(array_obj_ref_712_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_712_gather_scatter:flowthrough  inputs: " & " slice_714_wire = "& Convert_SLV_To_Hex_String(slice_714_wire) & "outputs: " & " array_obj_ref_712_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_712_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_712_gather_scatter
    process(slice_714_wire) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := slice_714_wire;
      ov(15 downto 0) := iv;
      array_obj_ref_712_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_717_gather_scatter flow-through 
    process(array_obj_ref_717_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_717_gather_scatter:flowthrough  inputs: " & " slice_719_wire = "& Convert_SLV_To_Hex_String(slice_719_wire) & "outputs: " & " array_obj_ref_717_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_717_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_717_gather_scatter
    process(slice_719_wire) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := slice_719_wire;
      ov(15 downto 0) := iv;
      array_obj_ref_717_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_722_gather_scatter flow-through 
    process(array_obj_ref_722_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_722_gather_scatter:flowthrough  inputs: " & " slice_724_wire = "& Convert_SLV_To_Hex_String(slice_724_wire) & "outputs: " & " array_obj_ref_722_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_722_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_722_gather_scatter
    process(slice_724_wire) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := slice_724_wire;
      ov(15 downto 0) := iv;
      array_obj_ref_722_data_0 <= ov(15 downto 0);
      --
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_344_branch_req_0," req0 do_while_stmt_344_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_344_branch_ack_0," ack0 do_while_stmt_344_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_344_branch_ack_1," ack1 do_while_stmt_344_branch");
    do_while_stmt_344_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u12_u1_441_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_344_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_344_branch_req_0,
          ack0 => do_while_stmt_344_branch_ack_0,
          ack1 => do_while_stmt_344_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_455_branch_req_0," req0 do_while_stmt_455_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_455_branch_ack_0," ack0 do_while_stmt_455_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_455_branch_ack_1," ack1 do_while_stmt_455_branch");
    do_while_stmt_455_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u12_u1_563_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_455_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_455_branch_req_0,
          ack0 => do_while_stmt_455_branch_ack_0,
          ack1 => do_while_stmt_455_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_577_branch_req_0," req0 do_while_stmt_577_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_577_branch_ack_0," ack0 do_while_stmt_577_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_577_branch_ack_1," ack1 do_while_stmt_577_branch");
    do_while_stmt_577_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u32_u1_616_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_577_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_577_branch_req_0,
          ack0 => do_while_stmt_577_branch_ack_0,
          ack1 => do_while_stmt_577_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_640_branch_req_0," req0 do_while_stmt_640_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_640_branch_ack_0," ack0 do_while_stmt_640_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_640_branch_ack_1," ack1 do_while_stmt_640_branch");
    do_while_stmt_640_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u12_u1_695_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_640_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_640_branch_req_0,
          ack0 => do_while_stmt_640_branch_ack_0,
          ack1 => do_while_stmt_640_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_731_branch_req_0," req0 if_stmt_731_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_731_branch_ack_0," ack0 if_stmt_731_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_731_branch_ack_1," ack1 if_stmt_731_branch");
    if_stmt_731_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u12_u1_734_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_731_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_731_branch_req_0,
          ack0 => if_stmt_731_branch_ack_0,
          ack1 => if_stmt_731_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_743_branch_req_0," req0 if_stmt_743_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_743_branch_ack_0," ack0 if_stmt_743_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_743_branch_ack_1," ack1 if_stmt_743_branch");
    if_stmt_743_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u12_u1_746_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_743_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_743_branch_req_0,
          ack0 => if_stmt_743_branch_ack_0,
          ack1 => if_stmt_743_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator ADD_u12_u12_358_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_358_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_358_inst:started:   inputs: " & " T_310_delayed_4_0_354 = "& Convert_SLV_To_Hex_String(T_310_delayed_4_0_354) & " LOAD_ZJ_357_wire = "& Convert_SLV_To_Hex_String(LOAD_ZJ_357_wire));
          --
        end if; 
        if ADD_u12_u12_358_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_358_inst:finished:  outputs: " & " NNNT_359= "  & Convert_SLV_To_Hex_String(NNNT_359));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (0) : ADD_u12_u12_358_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(23 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= T_310_delayed_4_0_354 & LOAD_ZJ_357_wire;
      NNNT_359 <= data_out(11 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u12_u12_358_inst_req_0;
      ADD_u12_u12_358_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_358_inst_req_1;
      ADD_u12_u12_358_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 12, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- logger for split-operator ADD_u12_u12_385_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_385_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_385_inst:started:   inputs: " & " T_346 = "& Convert_SLV_To_Hex_String(T_346) & " konst_384_wire_constant = "& Convert_SLV_To_Hex_String(konst_384_wire_constant));
          --
        end if; 
        if ADD_u12_u12_385_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_385_inst:finished:  outputs: " & " TT_386= "  & Convert_SLV_To_Hex_String(TT_386));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (1) : ADD_u12_u12_385_inst 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= T_346;
      TT_386 <= data_out(11 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u12_u12_385_inst_req_0;
      ADD_u12_u12_385_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_385_inst_req_1;
      ADD_u12_u12_385_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000000000001",
          constant_width => 12,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- logger for split-operator ADD_u12_u12_412_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_412_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_412_inst:started:   inputs: " & " T_346 = "& Convert_SLV_To_Hex_String(T_346) & " konst_411_wire_constant = "& Convert_SLV_To_Hex_String(konst_411_wire_constant));
          --
        end if; 
        if ADD_u12_u12_412_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_412_inst:finished:  outputs: " & " TTT_413= "  & Convert_SLV_To_Hex_String(TTT_413));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (2) : ADD_u12_u12_412_inst 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= T_346;
      TTT_413 <= data_out(11 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u12_u12_412_inst_req_0;
      ADD_u12_u12_412_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_412_inst_req_1;
      ADD_u12_u12_412_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_2_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000000000010",
          constant_width => 12,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- logger for split-operator ADD_u12_u12_417_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_417_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_417_inst:started:   inputs: " & " T_346 = "& Convert_SLV_To_Hex_String(T_346) & " konst_416_wire_constant = "& Convert_SLV_To_Hex_String(konst_416_wire_constant));
          --
        end if; 
        if ADD_u12_u12_417_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_417_inst:finished:  outputs: " & " TTTT_418= "  & Convert_SLV_To_Hex_String(TTTT_418));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (3) : ADD_u12_u12_417_inst 
    ApIntAdd_group_3: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= T_346;
      TTTT_418 <= data_out(11 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u12_u12_417_inst_req_0;
      ADD_u12_u12_417_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_417_inst_req_1;
      ADD_u12_u12_417_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_3_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000000000011",
          constant_width => 12,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- logger for split-operator ADD_u12_u12_436_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_436_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_436_inst:started:   inputs: " & " T_346 = "& Convert_SLV_To_Hex_String(T_346) & " konst_435_wire_constant = "& Convert_SLV_To_Hex_String(konst_435_wire_constant));
          --
        end if; 
        if ADD_u12_u12_436_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_436_inst:finished:  outputs: " & " NT_437= "  & Convert_SLV_To_Hex_String(NT_437));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (4) : ADD_u12_u12_436_inst 
    ApIntAdd_group_4: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= T_346;
      NT_437 <= data_out(11 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u12_u12_436_inst_req_0;
      ADD_u12_u12_436_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_436_inst_req_1;
      ADD_u12_u12_436_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_4_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000000000100",
          constant_width => 12,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- logger for split-operator ADD_u12_u12_553_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_553_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_553_inst:started:   inputs: " & " J_457 = "& Convert_SLV_To_Hex_String(J_457) & " konst_552_wire_constant = "& Convert_SLV_To_Hex_String(konst_552_wire_constant));
          --
        end if; 
        if ADD_u12_u12_553_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_553_inst:finished:  outputs: " & " NJ_554= "  & Convert_SLV_To_Hex_String(NJ_554));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (5) : ADD_u12_u12_553_inst 
    ApIntAdd_group_5: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= J_457;
      NJ_554 <= data_out(11 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u12_u12_553_inst_req_0;
      ADD_u12_u12_553_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_553_inst_req_1;
      ADD_u12_u12_553_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_5_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000000100000",
          constant_width => 12,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- logger for split-operator ADD_u12_u12_621_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_621_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_621_inst:started:   inputs: " & " L_567 = "& Convert_SLV_To_Hex_String(L_567) & " G_445 = "& Convert_SLV_To_Hex_String(G_445));
          --
        end if; 
        if ADD_u12_u12_621_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_621_inst:finished:  outputs: " & " ADD_u12_u12_621_wire= "  & Convert_SLV_To_Hex_String(ADD_u12_u12_621_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (6) : ADD_u12_u12_621_inst 
    ApIntAdd_group_6: Block -- 
      signal data_in: std_logic_vector(23 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= L_567 & G_445;
      ADD_u12_u12_621_wire <= data_out(11 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u12_u12_621_inst_req_0;
      ADD_u12_u12_621_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_621_inst_req_1;
      ADD_u12_u12_621_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_6_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 12, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- logger for split-operator ADD_u12_u12_629_inst flow-through 
    process(ADD_u12_u12_629_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_629_inst:flowthrough inputs: " & " L_567 = "& Convert_SLV_To_Hex_String(L_567) & " G_445 = "& Convert_SLV_To_Hex_String(G_445) & " outputs:" & " ADD_u12_u12_629_wire= "  & Convert_SLV_To_Hex_String(ADD_u12_u12_629_wire));
      --
    end process; 
    -- binary operator ADD_u12_u12_629_inst
    process(L_567, G_445) -- 
      variable tmp_var : std_logic_vector(11 downto 0); -- 
    begin -- 
      ApIntAdd_proc(L_567, G_445, tmp_var);
      ADD_u12_u12_629_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u12_u12_651_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_651_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_651_inst:started:   inputs: " & " H_642 = "& Convert_SLV_To_Hex_String(H_642) & " konst_650_wire_constant = "& Convert_SLV_To_Hex_String(konst_650_wire_constant));
          --
        end if; 
        if ADD_u12_u12_651_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_651_inst:finished:  outputs: " & " HH_652= "  & Convert_SLV_To_Hex_String(HH_652));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (8) : ADD_u12_u12_651_inst 
    ApIntAdd_group_8: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= H_642;
      HH_652 <= data_out(11 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u12_u12_651_inst_req_0;
      ADD_u12_u12_651_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_651_inst_req_1;
      ADD_u12_u12_651_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_8_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_8",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000000000001",
          constant_width => 12,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- logger for split-operator ADD_u12_u12_664_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_664_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_664_inst:started:   inputs: " & " H_642 = "& Convert_SLV_To_Hex_String(H_642) & " konst_663_wire_constant = "& Convert_SLV_To_Hex_String(konst_663_wire_constant));
          --
        end if; 
        if ADD_u12_u12_664_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_664_inst:finished:  outputs: " & " HHH_665= "  & Convert_SLV_To_Hex_String(HHH_665));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (9) : ADD_u12_u12_664_inst 
    ApIntAdd_group_9: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= H_642;
      HHH_665 <= data_out(11 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u12_u12_664_inst_req_0;
      ADD_u12_u12_664_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_664_inst_req_1;
      ADD_u12_u12_664_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_9_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_9",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000000000010",
          constant_width => 12,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- logger for split-operator ADD_u12_u12_677_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_677_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_677_inst:started:   inputs: " & " H_642 = "& Convert_SLV_To_Hex_String(H_642) & " konst_676_wire_constant = "& Convert_SLV_To_Hex_String(konst_676_wire_constant));
          --
        end if; 
        if ADD_u12_u12_677_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_677_inst:finished:  outputs: " & " HHHH_678= "  & Convert_SLV_To_Hex_String(HHHH_678));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (10) : ADD_u12_u12_677_inst 
    ApIntAdd_group_10: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= H_642;
      HHHH_678 <= data_out(11 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u12_u12_677_inst_req_0;
      ADD_u12_u12_677_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_677_inst_req_1;
      ADD_u12_u12_677_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_10_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_10",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000000000011",
          constant_width => 12,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- logger for split-operator ADD_u12_u12_690_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_690_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_690_inst:started:   inputs: " & " H_642 = "& Convert_SLV_To_Hex_String(H_642) & " konst_689_wire_constant = "& Convert_SLV_To_Hex_String(konst_689_wire_constant));
          --
        end if; 
        if ADD_u12_u12_690_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_690_inst:finished:  outputs: " & " NH_691= "  & Convert_SLV_To_Hex_String(NH_691));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (11) : ADD_u12_u12_690_inst 
    ApIntAdd_group_11: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= H_642;
      NH_691 <= data_out(11 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u12_u12_690_inst_req_0;
      ADD_u12_u12_690_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_690_inst_req_1;
      ADD_u12_u12_690_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_11_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_11",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000000000100",
          constant_width => 12,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- logger for split-operator ADD_u12_u12_700_inst flow-through 
    process(ADD_u12_u12_700_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_700_inst:flowthrough inputs: " & " L_567 = "& Convert_SLV_To_Hex_String(L_567) & " G_445 = "& Convert_SLV_To_Hex_String(G_445) & " outputs:" & " ADD_u12_u12_700_wire= "  & Convert_SLV_To_Hex_String(ADD_u12_u12_700_wire));
      --
    end process; 
    -- binary operator ADD_u12_u12_700_inst
    process(L_567, G_445) -- 
      variable tmp_var : std_logic_vector(11 downto 0); -- 
    begin -- 
      ApIntAdd_proc(L_567, G_445, tmp_var);
      ADD_u12_u12_700_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u12_u12_702_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_702_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_702_inst:started:   inputs: " & " ADD_u12_u12_700_wire = "& Convert_SLV_To_Hex_String(ADD_u12_u12_700_wire) & " konst_701_wire_constant = "& Convert_SLV_To_Hex_String(konst_701_wire_constant));
          --
        end if; 
        if ADD_u12_u12_702_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_702_inst:finished:  outputs: " & " ADD_u12_u12_702_wire= "  & Convert_SLV_To_Hex_String(ADD_u12_u12_702_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (13) : ADD_u12_u12_702_inst 
    ApIntAdd_group_13: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u12_u12_700_wire;
      ADD_u12_u12_702_wire <= data_out(11 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u12_u12_702_inst_req_0;
      ADD_u12_u12_702_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_702_inst_req_1;
      ADD_u12_u12_702_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_13_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000000000100",
          constant_width => 12,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- logger for split-operator ADD_u12_u12_729_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_729_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_729_inst:started:   inputs: " & " L_567 = "& Convert_SLV_To_Hex_String(L_567) & " konst_728_wire_constant = "& Convert_SLV_To_Hex_String(konst_728_wire_constant));
          --
        end if; 
        if ADD_u12_u12_729_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_729_inst:finished:  outputs: " & " NL_730= "  & Convert_SLV_To_Hex_String(NL_730));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (14) : ADD_u12_u12_729_inst 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= L_567;
      NL_730 <= data_out(11 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u12_u12_729_inst_req_0;
      ADD_u12_u12_729_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_729_inst_req_1;
      ADD_u12_u12_729_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_14_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000000000001",
          constant_width => 12,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- logger for split-operator ADD_u12_u12_741_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u12_u12_741_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_741_inst:started:   inputs: " & " G_445 = "& Convert_SLV_To_Hex_String(G_445) & " konst_740_wire_constant = "& Convert_SLV_To_Hex_String(konst_740_wire_constant));
          --
        end if; 
        if ADD_u12_u12_741_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u12_u12_741_inst:finished:  outputs: " & " NG_742= "  & Convert_SLV_To_Hex_String(NG_742));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (15) : ADD_u12_u12_741_inst 
    ApIntAdd_group_15: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= G_445;
      NG_742 <= data_out(11 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u12_u12_741_inst_req_0;
      ADD_u12_u12_741_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u12_u12_741_inst_req_1;
      ADD_u12_u12_741_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_15_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_15_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_15",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 12,
          constant_operand => "000000100000",
          constant_width => 12,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- logger for split-operator ADD_u16_u16_502_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u16_u16_502_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u16_u16_502_inst:started:   inputs: " & " LOAD_PJ_500_wire = "& Convert_SLV_To_Hex_String(LOAD_PJ_500_wire) & " konst_501_wire_constant = "& Convert_SLV_To_Hex_String(konst_501_wire_constant));
          --
        end if; 
        if ADD_u16_u16_502_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u16_u16_502_inst:finished:  outputs: " & " PPJ_503= "  & Convert_SLV_To_Hex_String(PPJ_503));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (16) : ADD_u16_u16_502_inst 
    ApIntAdd_group_16: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LOAD_PJ_500_wire;
      PPJ_503 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_502_inst_req_0;
      ADD_u16_u16_502_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_502_inst_req_1;
      ADD_u16_u16_502_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_16_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_16_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_16",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- logger for split-operator ADD_u16_u16_529_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u16_u16_529_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u16_u16_529_inst:started:   inputs: " & " LOAD_PJ_527_wire = "& Convert_SLV_To_Hex_String(LOAD_PJ_527_wire) & " konst_528_wire_constant = "& Convert_SLV_To_Hex_String(konst_528_wire_constant));
          --
        end if; 
        if ADD_u16_u16_529_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u16_u16_529_inst:finished:  outputs: " & " PPPJ_530= "  & Convert_SLV_To_Hex_String(PPPJ_530));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (17) : ADD_u16_u16_529_inst 
    ApIntAdd_group_17: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LOAD_PJ_527_wire;
      PPPJ_530 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_529_inst_req_0;
      ADD_u16_u16_529_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_529_inst_req_1;
      ADD_u16_u16_529_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_17_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_17_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_17",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- logger for split-operator ADD_u16_u16_534_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u16_u16_534_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u16_u16_534_inst:started:   inputs: " & " LOAD_PJ_532_wire = "& Convert_SLV_To_Hex_String(LOAD_PJ_532_wire) & " konst_533_wire_constant = "& Convert_SLV_To_Hex_String(konst_533_wire_constant));
          --
        end if; 
        if ADD_u16_u16_534_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u16_u16_534_inst:finished:  outputs: " & " PPPPJ_535= "  & Convert_SLV_To_Hex_String(PPPPJ_535));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (18) : ADD_u16_u16_534_inst 
    ApIntAdd_group_18: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LOAD_PJ_532_wire;
      PPPPJ_535 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_534_inst_req_0;
      ADD_u16_u16_534_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_534_inst_req_1;
      ADD_u16_u16_534_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_18_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_18_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_18",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- logger for split-operator ADD_u16_u16_558_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u16_u16_558_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u16_u16_558_inst:started:   inputs: " & " LOAD_PJ_556_wire = "& Convert_SLV_To_Hex_String(LOAD_PJ_556_wire) & " konst_557_wire_constant = "& Convert_SLV_To_Hex_String(konst_557_wire_constant));
          --
        end if; 
        if ADD_u16_u16_558_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u16_u16_558_inst:finished:  outputs: " & " ADD_u16_u16_558_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_558_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (19) : ADD_u16_u16_558_inst 
    ApIntAdd_group_19: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LOAD_PJ_556_wire;
      ADD_u16_u16_558_wire <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_558_inst_req_0;
      ADD_u16_u16_558_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_558_inst_req_1;
      ADD_u16_u16_558_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_19_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_19_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_19",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000100",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- logger for split-operator ADD_u16_u16_606_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u16_u16_606_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u16_u16_606_inst:started:   inputs: " & " LOAD_total_603_wire = "& Convert_SLV_To_Hex_String(LOAD_total_603_wire) & " array_obj_ref_605_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_605_wire));
          --
        end if; 
        if ADD_u16_u16_606_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u16_u16_606_inst:finished:  outputs: " & " ADD_u16_u16_606_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_606_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (20) : ADD_u16_u16_606_inst 
    ApIntAdd_group_20: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LOAD_total_603_wire & array_obj_ref_605_wire;
      ADD_u16_u16_606_wire <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u16_u16_606_inst_req_0;
      ADD_u16_u16_606_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u16_u16_606_inst_req_1;
      ADD_u16_u16_606_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_20_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_20_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_20",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- logger for split-operator ADD_u32_u32_485_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u32_u32_485_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u32_u32_485_inst:started:   inputs: " & " NNG_478 = "& Convert_SLV_To_Hex_String(NNG_478) & " NGG_420_delayed_4_0_481 = "& Convert_SLV_To_Hex_String(NGG_420_delayed_4_0_481));
          --
        end if; 
        if ADD_u32_u32_485_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u32_u32_485_inst:finished:  outputs: " & " NNJ_486= "  & Convert_SLV_To_Hex_String(NNJ_486));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (21) : ADD_u32_u32_485_inst 
    ApIntAdd_group_21: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= NNG_478 & NGG_420_delayed_4_0_481;
      NNJ_486 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_485_inst_req_0;
      ADD_u32_u32_485_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_485_inst_req_1;
      ADD_u32_u32_485_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_21_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_21_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_21",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- logger for split-operator ADD_u32_u32_611_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u32_u32_611_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u32_u32_611_inst:started:   inputs: " & " K_579 = "& Convert_SLV_To_Hex_String(K_579) & " konst_610_wire_constant = "& Convert_SLV_To_Hex_String(konst_610_wire_constant));
          --
        end if; 
        if ADD_u32_u32_611_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ADD_u32_u32_611_inst:finished:  outputs: " & " NK_612= "  & Convert_SLV_To_Hex_String(NK_612));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (22) : ADD_u32_u32_611_inst 
    ApIntAdd_group_22: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= K_579;
      NK_612 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_611_inst_req_0;
      ADD_u32_u32_611_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_611_inst_req_1;
      ADD_u32_u32_611_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_22_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_22_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_22",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- logger for split-operator CONCAT_u1_u32_368_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if CONCAT_u1_u32_368_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:CONCAT_u1_u32_368_inst:started:   inputs: " & " LOAD_one_366_wire = "& Convert_SLV_To_Hex_String(LOAD_one_366_wire) & " NTT_364 = "& Convert_SLV_To_Hex_String(NTT_364));
          --
        end if; 
        if CONCAT_u1_u32_368_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:CONCAT_u1_u32_368_inst:finished:  outputs: " & " NNT_369= "  & Convert_SLV_To_Hex_String(NNT_369));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (23) : CONCAT_u1_u32_368_inst 
    ApConcat_group_23: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LOAD_one_366_wire & NTT_364;
      NNT_369 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u1_u32_368_inst_req_0;
      CONCAT_u1_u32_368_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u1_u32_368_inst_req_1;
      CONCAT_u1_u32_368_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_23_gI: SplitGuardInterface generic map(name => "ApConcat_group_23_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_23",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 31, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- logger for split-operator CONCAT_u1_u32_477_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if CONCAT_u1_u32_477_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:CONCAT_u1_u32_477_inst:started:   inputs: " & " LOAD_one_475_wire = "& Convert_SLV_To_Hex_String(LOAD_one_475_wire) & " NJJ_415_delayed_2_0_473 = "& Convert_SLV_To_Hex_String(NJJ_415_delayed_2_0_473));
          --
        end if; 
        if CONCAT_u1_u32_477_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:CONCAT_u1_u32_477_inst:finished:  outputs: " & " NNG_478= "  & Convert_SLV_To_Hex_String(NNG_478));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (24) : CONCAT_u1_u32_477_inst 
    ApConcat_group_24: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LOAD_one_475_wire & NJJ_415_delayed_2_0_473;
      NNG_478 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u1_u32_477_inst_req_0;
      CONCAT_u1_u32_477_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u1_u32_477_inst_req_1;
      CONCAT_u1_u32_477_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_24_gI: SplitGuardInterface generic map(name => "ApConcat_group_24_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_24",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 31, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- logger for split-operator CONCAT_u4_u16_630_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if CONCAT_u4_u16_630_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:CONCAT_u4_u16_630_inst:started:   inputs: " & " LOAD_zer_626_wire = "& Convert_SLV_To_Hex_String(LOAD_zer_626_wire) & " ADD_u12_u12_629_wire = "& Convert_SLV_To_Hex_String(ADD_u12_u12_629_wire));
          --
        end if; 
        if CONCAT_u4_u16_630_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:CONCAT_u4_u16_630_inst:finished:  outputs: " & " f_631= "  & Convert_SLV_To_Hex_String(f_631));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (25) : CONCAT_u4_u16_630_inst 
    ApConcat_group_25: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LOAD_zer_626_wire & ADD_u12_u12_629_wire;
      f_631 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u4_u16_630_inst_req_0;
      CONCAT_u4_u16_630_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u4_u16_630_inst_req_1;
      CONCAT_u4_u16_630_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_25_gI: SplitGuardInterface generic map(name => "ApConcat_group_25_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_25",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 12, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- logger for split-operator MUL_u16_u16_600_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if MUL_u16_u16_600_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:MUL_u16_u16_600_inst:started:   inputs: " & " imag1_588 = "& Convert_SLV_To_Hex_String(imag1_588) & " ker1_592 = "& Convert_SLV_To_Hex_String(ker1_592));
          --
        end if; 
        if MUL_u16_u16_600_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:MUL_u16_u16_600_inst:finished:  outputs: " & " MUL_u16_u16_600_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_600_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (26) : MUL_u16_u16_600_inst 
    ApIntMul_group_26: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= imag1_588 & ker1_592;
      MUL_u16_u16_600_wire <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= MUL_u16_u16_600_inst_req_0;
      MUL_u16_u16_600_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= MUL_u16_u16_600_inst_req_1;
      MUL_u16_u16_600_inst_ack_1 <= ackR_unguarded(0);
      ApIntMul_group_26_gI: SplitGuardInterface generic map(name => "ApIntMul_group_26_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          name => "ApIntMul_group_26",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- logger for split-operator ULT_u12_u1_441_inst flow-through 
    process(ULT_u12_u1_441_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ULT_u12_u1_441_inst:flowthrough inputs: " & " NT_437 = "& Convert_SLV_To_Hex_String(NT_437) & " konst_440_wire_constant = "& Convert_SLV_To_Hex_String(konst_440_wire_constant) & " outputs:" & " ULT_u12_u1_441_wire= "  & Convert_SLV_To_Hex_String(ULT_u12_u1_441_wire));
      --
    end process; 
    -- binary operator ULT_u12_u1_441_inst
    process(NT_437) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(NT_437, konst_440_wire_constant, tmp_var);
      ULT_u12_u1_441_wire <= tmp_var; --
    end process;
    -- logger for split-operator ULT_u12_u1_563_inst flow-through 
    process(ULT_u12_u1_563_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ULT_u12_u1_563_inst:flowthrough inputs: " & " NJ_554 = "& Convert_SLV_To_Hex_String(NJ_554) & " konst_562_wire_constant = "& Convert_SLV_To_Hex_String(konst_562_wire_constant) & " outputs:" & " ULT_u12_u1_563_wire= "  & Convert_SLV_To_Hex_String(ULT_u12_u1_563_wire));
      --
    end process; 
    -- binary operator ULT_u12_u1_563_inst
    process(NJ_554) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(NJ_554, konst_562_wire_constant, tmp_var);
      ULT_u12_u1_563_wire <= tmp_var; --
    end process;
    -- logger for split-operator ULT_u12_u1_695_inst flow-through 
    process(ULT_u12_u1_695_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ULT_u12_u1_695_inst:flowthrough inputs: " & " NH_691 = "& Convert_SLV_To_Hex_String(NH_691) & " konst_694_wire_constant = "& Convert_SLV_To_Hex_String(konst_694_wire_constant) & " outputs:" & " ULT_u12_u1_695_wire= "  & Convert_SLV_To_Hex_String(ULT_u12_u1_695_wire));
      --
    end process; 
    -- binary operator ULT_u12_u1_695_inst
    process(NH_691) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(NH_691, konst_694_wire_constant, tmp_var);
      ULT_u12_u1_695_wire <= tmp_var; --
    end process;
    -- logger for split-operator ULT_u12_u1_734_inst flow-through 
    process(ULT_u12_u1_734_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ULT_u12_u1_734_inst:flowthrough inputs: " & " NL_730 = "& Convert_SLV_To_Hex_String(NL_730) & " konst_733_wire_constant = "& Convert_SLV_To_Hex_String(konst_733_wire_constant) & " outputs:" & " ULT_u12_u1_734_wire= "  & Convert_SLV_To_Hex_String(ULT_u12_u1_734_wire));
      --
    end process; 
    -- binary operator ULT_u12_u1_734_inst
    process(NL_730) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(NL_730, konst_733_wire_constant, tmp_var);
      ULT_u12_u1_734_wire <= tmp_var; --
    end process;
    -- logger for split-operator ULT_u12_u1_746_inst flow-through 
    process(ULT_u12_u1_746_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ULT_u12_u1_746_inst:flowthrough inputs: " & " NG_742 = "& Convert_SLV_To_Hex_String(NG_742) & " konst_745_wire_constant = "& Convert_SLV_To_Hex_String(konst_745_wire_constant) & " outputs:" & " ULT_u12_u1_746_wire= "  & Convert_SLV_To_Hex_String(ULT_u12_u1_746_wire));
      --
    end process; 
    -- binary operator ULT_u12_u1_746_inst
    process(NG_742) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(NG_742, konst_745_wire_constant, tmp_var);
      ULT_u12_u1_746_wire <= tmp_var; --
    end process;
    -- logger for split-operator ULT_u32_u1_616_inst flow-through 
    process(ULT_u32_u1_616_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:ULT_u32_u1_616_inst:flowthrough inputs: " & " NK_612 = "& Convert_SLV_To_Hex_String(NK_612) & " konst_615_wire_constant = "& Convert_SLV_To_Hex_String(konst_615_wire_constant) & " outputs:" & " ULT_u32_u1_616_wire= "  & Convert_SLV_To_Hex_String(ULT_u32_u1_616_wire));
      --
    end process; 
    -- binary operator ULT_u32_u1_616_inst
    process(NK_612) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(NK_612, konst_615_wire_constant, tmp_var);
      ULT_u32_u1_616_wire <= tmp_var; --
    end process;
    -- logger for split-operator LOAD_PJ_527_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if LOAD_PJ_527_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_PJ_527_load_0:started:   inputs: " & " LOAD_PJ_527_word_address_0 = "& Convert_SLV_To_Hex_String(LOAD_PJ_527_word_address_0));
          --
        end if; 
        if LOAD_PJ_527_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_PJ_527_load_0:finished:  outputs: " & " LOAD_PJ_527_data_0= "  & Convert_SLV_To_Hex_String(LOAD_PJ_527_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator LOAD_PJ_532_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if LOAD_PJ_532_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_PJ_532_load_0:started:   inputs: " & " LOAD_PJ_532_word_address_0 = "& Convert_SLV_To_Hex_String(LOAD_PJ_532_word_address_0));
          --
        end if; 
        if LOAD_PJ_532_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_PJ_532_load_0:finished:  outputs: " & " LOAD_PJ_532_data_0= "  & Convert_SLV_To_Hex_String(LOAD_PJ_532_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator LOAD_PJ_556_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if LOAD_PJ_556_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_PJ_556_load_0:started:   inputs: " & " LOAD_PJ_556_word_address_0 = "& Convert_SLV_To_Hex_String(LOAD_PJ_556_word_address_0));
          --
        end if; 
        if LOAD_PJ_556_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_PJ_556_load_0:finished:  outputs: " & " LOAD_PJ_556_data_0= "  & Convert_SLV_To_Hex_String(LOAD_PJ_556_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator LOAD_PJ_500_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if LOAD_PJ_500_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_PJ_500_load_0:started:   inputs: " & " LOAD_PJ_500_word_address_0 = "& Convert_SLV_To_Hex_String(LOAD_PJ_500_word_address_0));
          --
        end if; 
        if LOAD_PJ_500_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_PJ_500_load_0:finished:  outputs: " & " LOAD_PJ_500_data_0= "  & Convert_SLV_To_Hex_String(LOAD_PJ_500_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator LOAD_PJ_505_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if LOAD_PJ_505_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_PJ_505_load_0:started:   inputs: " & " LOAD_PJ_505_word_address_0 = "& Convert_SLV_To_Hex_String(LOAD_PJ_505_word_address_0));
          --
        end if; 
        if LOAD_PJ_505_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_PJ_505_load_0:finished:  outputs: " & " LOAD_PJ_505_data_0= "  & Convert_SLV_To_Hex_String(LOAD_PJ_505_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (0) : LOAD_PJ_527_load_0 LOAD_PJ_532_load_0 LOAD_PJ_556_load_0 LOAD_PJ_500_load_0 LOAD_PJ_505_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(4 downto 0);
      signal data_out: std_logic_vector(79 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 4 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 4 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 4 downto 0);
      signal guard_vector : std_logic_vector( 4 downto 0);
      constant inBUFs : IntegerArray(4 downto 0) := (4 => 2, 3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(4 downto 0) := (4 => 2, 3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(4 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false);
      constant guardBuffering: IntegerArray(4 downto 0)  := (0 => 4, 1 => 4, 2 => 4, 3 => 4, 4 => 4);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        LOAD_PJ_527_load_0_req_0,
        LOAD_PJ_527_load_0_ack_0,
        LOAD_PJ_527_load_0_req_1,
        LOAD_PJ_527_load_0_ack_1,
        "LOAD_PJ_527_load_0",
        "memory_space_0" ,
        LOAD_PJ_527_data_0,
        LOAD_PJ_527_word_address_0,
        "LOAD_PJ_527_data_0",
        "LOAD_PJ_527_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        LOAD_PJ_532_load_0_req_0,
        LOAD_PJ_532_load_0_ack_0,
        LOAD_PJ_532_load_0_req_1,
        LOAD_PJ_532_load_0_ack_1,
        "LOAD_PJ_532_load_0",
        "memory_space_0" ,
        LOAD_PJ_532_data_0,
        LOAD_PJ_532_word_address_0,
        "LOAD_PJ_532_data_0",
        "LOAD_PJ_532_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        LOAD_PJ_556_load_0_req_0,
        LOAD_PJ_556_load_0_ack_0,
        LOAD_PJ_556_load_0_req_1,
        LOAD_PJ_556_load_0_ack_1,
        "LOAD_PJ_556_load_0",
        "memory_space_0" ,
        LOAD_PJ_556_data_0,
        LOAD_PJ_556_word_address_0,
        "LOAD_PJ_556_data_0",
        "LOAD_PJ_556_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        LOAD_PJ_500_load_0_req_0,
        LOAD_PJ_500_load_0_ack_0,
        LOAD_PJ_500_load_0_req_1,
        LOAD_PJ_500_load_0_ack_1,
        "LOAD_PJ_500_load_0",
        "memory_space_0" ,
        LOAD_PJ_500_data_0,
        LOAD_PJ_500_word_address_0,
        "LOAD_PJ_500_data_0",
        "LOAD_PJ_500_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        LOAD_PJ_505_load_0_req_0,
        LOAD_PJ_505_load_0_ack_0,
        LOAD_PJ_505_load_0_req_1,
        LOAD_PJ_505_load_0_ack_1,
        "LOAD_PJ_505_load_0",
        "memory_space_0" ,
        LOAD_PJ_505_data_0,
        LOAD_PJ_505_word_address_0,
        "LOAD_PJ_505_data_0",
        "LOAD_PJ_505_word_address_0" -- 
      );
      reqL_unguarded(4) <= LOAD_PJ_527_load_0_req_0;
      reqL_unguarded(3) <= LOAD_PJ_532_load_0_req_0;
      reqL_unguarded(2) <= LOAD_PJ_556_load_0_req_0;
      reqL_unguarded(1) <= LOAD_PJ_500_load_0_req_0;
      reqL_unguarded(0) <= LOAD_PJ_505_load_0_req_0;
      LOAD_PJ_527_load_0_ack_0 <= ackL_unguarded(4);
      LOAD_PJ_532_load_0_ack_0 <= ackL_unguarded(3);
      LOAD_PJ_556_load_0_ack_0 <= ackL_unguarded(2);
      LOAD_PJ_500_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_PJ_505_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(4) <= LOAD_PJ_527_load_0_req_1;
      reqR_unguarded(3) <= LOAD_PJ_532_load_0_req_1;
      reqR_unguarded(2) <= LOAD_PJ_556_load_0_req_1;
      reqR_unguarded(1) <= LOAD_PJ_500_load_0_req_1;
      reqR_unguarded(0) <= LOAD_PJ_505_load_0_req_1;
      LOAD_PJ_527_load_0_ack_1 <= ackR_unguarded(4);
      LOAD_PJ_532_load_0_ack_1 <= ackR_unguarded(3);
      LOAD_PJ_556_load_0_ack_1 <= ackR_unguarded(2);
      LOAD_PJ_500_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_PJ_505_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 2) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 2) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_4", num_slots => 2) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 5, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_PJ_527_word_address_0 & LOAD_PJ_532_word_address_0 & LOAD_PJ_556_word_address_0 & LOAD_PJ_500_word_address_0 & LOAD_PJ_505_word_address_0;
      LOAD_PJ_527_data_0 <= data_out(79 downto 64);
      LOAD_PJ_532_data_0 <= data_out(63 downto 48);
      LOAD_PJ_556_data_0 <= data_out(47 downto 32);
      LOAD_PJ_500_data_0 <= data_out(31 downto 16);
      LOAD_PJ_505_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 5,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 5,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(15 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logger for split-operator LOAD_ZJ_357_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if LOAD_ZJ_357_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_ZJ_357_load_0:started:   inputs: " & " LOAD_ZJ_357_word_address_0 = "& Convert_SLV_To_Hex_String(LOAD_ZJ_357_word_address_0));
          --
        end if; 
        if LOAD_ZJ_357_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_ZJ_357_load_0:finished:  outputs: " & " LOAD_ZJ_357_data_0= "  & Convert_SLV_To_Hex_String(LOAD_ZJ_357_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (1) : LOAD_ZJ_357_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(11 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        LOAD_ZJ_357_load_0_req_0,
        LOAD_ZJ_357_load_0_ack_0,
        LOAD_ZJ_357_load_0_req_1,
        LOAD_ZJ_357_load_0_ack_1,
        "LOAD_ZJ_357_load_0",
        "memory_space_1" ,
        LOAD_ZJ_357_data_0,
        LOAD_ZJ_357_word_address_0,
        "LOAD_ZJ_357_data_0",
        "LOAD_ZJ_357_word_address_0" -- 
      );
      reqL_unguarded(0) <= LOAD_ZJ_357_load_0_req_0;
      LOAD_ZJ_357_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_ZJ_357_load_0_req_1;
      LOAD_ZJ_357_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_ZJ_357_word_address_0;
      LOAD_ZJ_357_data_0 <= data_out(11 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 1,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(0 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 12,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(11 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- logger for split-operator LOAD_one_366_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if LOAD_one_366_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_one_366_load_0:started:   inputs: " & " LOAD_one_366_word_address_0 = "& Convert_SLV_To_Hex_String(LOAD_one_366_word_address_0));
          --
        end if; 
        if LOAD_one_366_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_one_366_load_0:finished:  outputs: " & " LOAD_one_366_data_0= "  & Convert_SLV_To_Hex_String(LOAD_one_366_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator LOAD_one_475_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if LOAD_one_475_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_one_475_load_0:started:   inputs: " & " LOAD_one_475_word_address_0 = "& Convert_SLV_To_Hex_String(LOAD_one_475_word_address_0));
          --
        end if; 
        if LOAD_one_475_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_one_475_load_0:finished:  outputs: " & " LOAD_one_475_data_0= "  & Convert_SLV_To_Hex_String(LOAD_one_475_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (2) : LOAD_one_366_load_0 LOAD_one_475_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 4, 1 => 4);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        LOAD_one_366_load_0_req_0,
        LOAD_one_366_load_0_ack_0,
        LOAD_one_366_load_0_req_1,
        LOAD_one_366_load_0_ack_1,
        "LOAD_one_366_load_0",
        "memory_space_6" ,
        LOAD_one_366_data_0,
        LOAD_one_366_word_address_0,
        "LOAD_one_366_data_0",
        "LOAD_one_366_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        LOAD_one_475_load_0_req_0,
        LOAD_one_475_load_0_ack_0,
        LOAD_one_475_load_0_req_1,
        LOAD_one_475_load_0_ack_1,
        "LOAD_one_475_load_0",
        "memory_space_6" ,
        LOAD_one_475_data_0,
        LOAD_one_475_word_address_0,
        "LOAD_one_475_data_0",
        "LOAD_one_475_word_address_0" -- 
      );
      reqL_unguarded(1) <= LOAD_one_366_load_0_req_0;
      reqL_unguarded(0) <= LOAD_one_475_load_0_req_0;
      LOAD_one_366_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_one_475_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= LOAD_one_366_load_0_req_1;
      reqR_unguarded(0) <= LOAD_one_475_load_0_req_1;
      LOAD_one_366_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_one_475_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_one_366_word_address_0 & LOAD_one_475_word_address_0;
      LOAD_one_366_data_0 <= data_out(1 downto 1);
      LOAD_one_475_data_0 <= data_out(0 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 1,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(0 downto 0),
          mtag => memory_space_6_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- logger for split-operator LOAD_total_622_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if LOAD_total_622_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_total_622_load_0:started:   inputs: " & " LOAD_total_622_word_address_0 = "& Convert_SLV_To_Hex_String(LOAD_total_622_word_address_0));
          --
        end if; 
        if LOAD_total_622_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_total_622_load_0:finished:  outputs: " & " LOAD_total_622_data_0= "  & Convert_SLV_To_Hex_String(LOAD_total_622_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator LOAD_total_603_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if LOAD_total_603_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_total_603_load_0:started:   inputs: " & " LOAD_total_603_word_address_0 = "& Convert_SLV_To_Hex_String(LOAD_total_603_word_address_0));
          --
        end if; 
        if LOAD_total_603_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_total_603_load_0:finished:  outputs: " & " LOAD_total_603_data_0= "  & Convert_SLV_To_Hex_String(LOAD_total_603_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (3) : LOAD_total_622_load_0 LOAD_total_603_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 4, 1 => 2);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        LOAD_total_622_load_0_req_0,
        LOAD_total_622_load_0_ack_0,
        LOAD_total_622_load_0_req_1,
        LOAD_total_622_load_0_ack_1,
        "LOAD_total_622_load_0",
        "memory_space_7" ,
        LOAD_total_622_data_0,
        LOAD_total_622_word_address_0,
        "LOAD_total_622_data_0",
        "LOAD_total_622_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        LOAD_total_603_load_0_req_0,
        LOAD_total_603_load_0_ack_0,
        LOAD_total_603_load_0_req_1,
        LOAD_total_603_load_0_ack_1,
        "LOAD_total_603_load_0",
        "memory_space_7" ,
        LOAD_total_603_data_0,
        LOAD_total_603_word_address_0,
        "LOAD_total_603_data_0",
        "LOAD_total_603_word_address_0" -- 
      );
      reqL_unguarded(1) <= LOAD_total_622_load_0_req_0;
      reqL_unguarded(0) <= LOAD_total_603_load_0_req_0;
      LOAD_total_622_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_total_603_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= LOAD_total_622_load_0_req_1;
      reqR_unguarded(0) <= LOAD_total_603_load_0_req_1;
      LOAD_total_622_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_total_603_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_total_622_word_address_0 & LOAD_total_603_word_address_0;
      LOAD_total_622_data_0 <= data_out(31 downto 16);
      LOAD_total_603_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- logger for split-operator LOAD_zer_626_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if LOAD_zer_626_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_zer_626_load_0:started:   inputs: " & " LOAD_zer_626_word_address_0 = "& Convert_SLV_To_Hex_String(LOAD_zer_626_word_address_0));
          --
        end if; 
        if LOAD_zer_626_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:LOAD_zer_626_load_0:finished:  outputs: " & " LOAD_zer_626_data_0= "  & Convert_SLV_To_Hex_String(LOAD_zer_626_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (4) : LOAD_zer_626_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        LOAD_zer_626_load_0_req_0,
        LOAD_zer_626_load_0_ack_0,
        LOAD_zer_626_load_0_req_1,
        LOAD_zer_626_load_0_ack_1,
        "LOAD_zer_626_load_0",
        "memory_space_8" ,
        LOAD_zer_626_data_0,
        LOAD_zer_626_word_address_0,
        "LOAD_zer_626_data_0",
        "LOAD_zer_626_word_address_0" -- 
      );
      reqL_unguarded(0) <= LOAD_zer_626_load_0_req_0;
      LOAD_zer_626_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_zer_626_load_0_req_1;
      LOAD_zer_626_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_zer_626_word_address_0;
      LOAD_zer_626_data_0 <= data_out(3 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 4,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(3 downto 0),
          mtag => memory_space_8_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- logger for split-operator array_obj_ref_587_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_587_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_587_load_0:started:   inputs: " & " array_obj_ref_587_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_587_word_address_0));
          --
        end if; 
        if array_obj_ref_587_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_587_load_0:finished:  outputs: " & " array_obj_ref_587_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_587_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_685_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_685_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_685_load_0:started:   inputs: " & " array_obj_ref_685_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_685_word_address_0));
          --
        end if; 
        if array_obj_ref_685_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_685_load_0:finished:  outputs: " & " array_obj_ref_685_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_685_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_672_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_672_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_672_load_0:started:   inputs: " & " array_obj_ref_672_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_672_word_address_0));
          --
        end if; 
        if array_obj_ref_672_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_672_load_0:finished:  outputs: " & " array_obj_ref_672_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_672_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_659_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_659_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_659_load_0:started:   inputs: " & " array_obj_ref_659_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_659_word_address_0));
          --
        end if; 
        if array_obj_ref_659_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_659_load_0:finished:  outputs: " & " array_obj_ref_659_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_659_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (5) : array_obj_ref_587_load_0 array_obj_ref_685_load_0 array_obj_ref_672_load_0 array_obj_ref_659_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 4, 1 => 4, 2 => 4, 3 => 4);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_587_load_0_req_0,
        array_obj_ref_587_load_0_ack_0,
        array_obj_ref_587_load_0_req_1,
        array_obj_ref_587_load_0_ack_1,
        "array_obj_ref_587_load_0",
        "memory_space_3" ,
        array_obj_ref_587_data_0,
        array_obj_ref_587_word_address_0,
        "array_obj_ref_587_data_0",
        "array_obj_ref_587_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_685_load_0_req_0,
        array_obj_ref_685_load_0_ack_0,
        array_obj_ref_685_load_0_req_1,
        array_obj_ref_685_load_0_ack_1,
        "array_obj_ref_685_load_0",
        "memory_space_3" ,
        array_obj_ref_685_data_0,
        array_obj_ref_685_word_address_0,
        "array_obj_ref_685_data_0",
        "array_obj_ref_685_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_672_load_0_req_0,
        array_obj_ref_672_load_0_ack_0,
        array_obj_ref_672_load_0_req_1,
        array_obj_ref_672_load_0_ack_1,
        "array_obj_ref_672_load_0",
        "memory_space_3" ,
        array_obj_ref_672_data_0,
        array_obj_ref_672_word_address_0,
        "array_obj_ref_672_data_0",
        "array_obj_ref_672_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_659_load_0_req_0,
        array_obj_ref_659_load_0_ack_0,
        array_obj_ref_659_load_0_req_1,
        array_obj_ref_659_load_0_ack_1,
        "array_obj_ref_659_load_0",
        "memory_space_3" ,
        array_obj_ref_659_data_0,
        array_obj_ref_659_word_address_0,
        "array_obj_ref_659_data_0",
        "array_obj_ref_659_word_address_0" -- 
      );
      reqL_unguarded(3) <= array_obj_ref_587_load_0_req_0;
      reqL_unguarded(2) <= array_obj_ref_685_load_0_req_0;
      reqL_unguarded(1) <= array_obj_ref_672_load_0_req_0;
      reqL_unguarded(0) <= array_obj_ref_659_load_0_req_0;
      array_obj_ref_587_load_0_ack_0 <= ackL_unguarded(3);
      array_obj_ref_685_load_0_ack_0 <= ackL_unguarded(2);
      array_obj_ref_672_load_0_ack_0 <= ackL_unguarded(1);
      array_obj_ref_659_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= array_obj_ref_587_load_0_req_1;
      reqR_unguarded(2) <= array_obj_ref_685_load_0_req_1;
      reqR_unguarded(1) <= array_obj_ref_672_load_0_req_1;
      reqR_unguarded(0) <= array_obj_ref_659_load_0_req_1;
      array_obj_ref_587_load_0_ack_1 <= ackR_unguarded(3);
      array_obj_ref_685_load_0_ack_1 <= ackR_unguarded(2);
      array_obj_ref_672_load_0_ack_1 <= ackR_unguarded(1);
      array_obj_ref_659_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup5_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_2", num_slots => 2) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_3", num_slots => 2) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_587_word_address_0 & array_obj_ref_685_word_address_0 & array_obj_ref_672_word_address_0 & array_obj_ref_659_word_address_0;
      array_obj_ref_587_data_0 <= data_out(63 downto 48);
      array_obj_ref_685_data_0 <= data_out(47 downto 32);
      array_obj_ref_672_data_0 <= data_out(31 downto 16);
      array_obj_ref_659_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 4,
        num_reqs => 4,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(3 downto 0),
          mtag => memory_space_3_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 16,
        num_reqs => 4,
        tag_length => 4,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(15 downto 0),
          mtag => memory_space_3_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- logger for split-operator array_obj_ref_591_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_591_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_591_load_0:started:   inputs: " & " array_obj_ref_591_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_591_word_address_0));
          --
        end if; 
        if array_obj_ref_591_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_591_load_0:finished:  outputs: " & " array_obj_ref_591_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_591_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (6) : array_obj_ref_591_load_0 
    LoadGroup6: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_591_load_0_req_0,
        array_obj_ref_591_load_0_ack_0,
        array_obj_ref_591_load_0_req_1,
        array_obj_ref_591_load_0_ack_1,
        "array_obj_ref_591_load_0",
        "memory_space_4" ,
        array_obj_ref_591_data_0,
        array_obj_ref_591_word_address_0,
        "array_obj_ref_591_data_0",
        "array_obj_ref_591_word_address_0" -- 
      );
      reqL_unguarded(0) <= array_obj_ref_591_load_0_req_0;
      array_obj_ref_591_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_591_load_0_req_1;
      array_obj_ref_591_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup6_gI: SplitGuardInterface generic map(name => "LoadGroup6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_591_word_address_0;
      array_obj_ref_591_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup6", addr_width => 4,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(3 downto 0),
          mtag => memory_space_4_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup6 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(15 downto 0),
          mtag => memory_space_4_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 6
    -- logger for split-operator array_obj_ref_605_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_605_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_605_load_0:started:   inputs: " & " array_obj_ref_605_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_605_word_address_0));
          --
        end if; 
        if array_obj_ref_605_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_605_load_0:finished:  outputs: " & " array_obj_ref_605_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_605_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (7) : array_obj_ref_605_load_0 
    LoadGroup7: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_605_load_0_req_0,
        array_obj_ref_605_load_0_ack_0,
        array_obj_ref_605_load_0_req_1,
        array_obj_ref_605_load_0_ack_1,
        "array_obj_ref_605_load_0",
        "memory_space_2" ,
        array_obj_ref_605_data_0,
        array_obj_ref_605_word_address_0,
        "array_obj_ref_605_data_0",
        "array_obj_ref_605_word_address_0" -- 
      );
      reqL_unguarded(0) <= array_obj_ref_605_load_0_req_0;
      array_obj_ref_605_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_605_load_0_req_1;
      array_obj_ref_605_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup7_gI: SplitGuardInterface generic map(name => "LoadGroup7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_605_word_address_0;
      array_obj_ref_605_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup7", addr_width => 4,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(3 downto 0),
          mtag => memory_space_2_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup7 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(15 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 7
    -- logger for split-operator array_obj_ref_637_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_637_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_637_load_0:started:   inputs: " & " array_obj_ref_637_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_637_word_address_0));
          --
        end if; 
        if array_obj_ref_637_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_637_load_0:finished:  outputs: " & " array_obj_ref_637_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_637_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (8) : array_obj_ref_637_load_0 
    LoadGroup8: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_637_load_0_req_0,
        array_obj_ref_637_load_0_ack_0,
        array_obj_ref_637_load_0_req_1,
        array_obj_ref_637_load_0_ack_1,
        "array_obj_ref_637_load_0",
        "memory_space_5" ,
        array_obj_ref_637_data_0,
        array_obj_ref_637_word_address_0,
        "array_obj_ref_637_data_0",
        "array_obj_ref_637_word_address_0" -- 
      );
      reqL_unguarded(0) <= array_obj_ref_637_load_0_req_0;
      array_obj_ref_637_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_637_load_0_req_1;
      array_obj_ref_637_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup8_gI: SplitGuardInterface generic map(name => "LoadGroup8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_637_word_address_0;
      array_obj_ref_637_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup8", addr_width => 11,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(10 downto 0),
          mtag => memory_space_5_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup8 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(15 downto 0),
          mtag => memory_space_5_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 8
    -- logger for split-operator STORE_PJ_555_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if STORE_PJ_555_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:STORE_PJ_555_store_0:started:   inputs: " & " STORE_PJ_555_word_address_0 = "& Convert_SLV_To_Hex_String(STORE_PJ_555_word_address_0) & " STORE_PJ_555_data_0 = "& Convert_SLV_To_Hex_String(STORE_PJ_555_data_0));
          --
        end if; 
        if STORE_PJ_555_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:STORE_PJ_555_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator STORE_PJ_451_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if STORE_PJ_451_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:STORE_PJ_451_store_0:started:   inputs: " & " STORE_PJ_451_word_address_0 = "& Convert_SLV_To_Hex_String(STORE_PJ_451_word_address_0) & " STORE_PJ_451_data_0 = "& Convert_SLV_To_Hex_String(STORE_PJ_451_data_0));
          --
        end if; 
        if STORE_PJ_451_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:STORE_PJ_451_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      STORE_PJ_555_store_0_req_0,
      STORE_PJ_555_store_0_ack_0,
      STORE_PJ_555_store_0_req_1,
      STORE_PJ_555_store_0_ack_1,
      "STORE_PJ_555_store_0",
      "memory_space_0" ,
      STORE_PJ_555_data_0,
      STORE_PJ_555_word_address_0,
      "STORE_PJ_555_data_0",
      "STORE_PJ_555_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      STORE_PJ_451_store_0_req_0,
      STORE_PJ_451_store_0_ack_0,
      STORE_PJ_451_store_0_req_1,
      STORE_PJ_451_store_0_ack_1,
      "STORE_PJ_451_store_0",
      "memory_space_0" ,
      STORE_PJ_451_data_0,
      STORE_PJ_451_word_address_0,
      "STORE_PJ_451_data_0",
      "STORE_PJ_451_word_address_0" -- 
    );
    -- shared store operator group (0) : STORE_PJ_555_store_0 STORE_PJ_451_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(1 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 7, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 4);
      -- 
    begin -- 
      reqL_unguarded(1) <= STORE_PJ_555_store_0_req_0;
      reqL_unguarded(0) <= STORE_PJ_451_store_0_req_0;
      STORE_PJ_555_store_0_ack_0 <= ackL_unguarded(1);
      STORE_PJ_451_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= STORE_PJ_555_store_0_req_1;
      reqR_unguarded(0) <= STORE_PJ_451_store_0_req_1;
      STORE_PJ_555_store_0_ack_1 <= ackR_unguarded(1);
      STORE_PJ_451_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_PJ_555_word_address_0 & STORE_PJ_451_word_address_0;
      data_in <= STORE_PJ_555_data_0 & STORE_PJ_451_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(0 downto 0),
          mdata => memory_space_0_sr_data(15 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- logger for split-operator STORE_total_602_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if STORE_total_602_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:STORE_total_602_store_0:started:   inputs: " & " STORE_total_602_word_address_0 = "& Convert_SLV_To_Hex_String(STORE_total_602_word_address_0) & " STORE_total_602_data_0 = "& Convert_SLV_To_Hex_String(STORE_total_602_data_0));
          --
        end if; 
        if STORE_total_602_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:STORE_total_602_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator STORE_total_573_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if STORE_total_573_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:STORE_total_573_store_0:started:   inputs: " & " STORE_total_573_word_address_0 = "& Convert_SLV_To_Hex_String(STORE_total_573_word_address_0) & " STORE_total_573_data_0 = "& Convert_SLV_To_Hex_String(STORE_total_573_data_0));
          --
        end if; 
        if STORE_total_573_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:STORE_total_573_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      STORE_total_602_store_0_req_0,
      STORE_total_602_store_0_ack_0,
      STORE_total_602_store_0_req_1,
      STORE_total_602_store_0_ack_1,
      "STORE_total_602_store_0",
      "memory_space_7" ,
      STORE_total_602_data_0,
      STORE_total_602_word_address_0,
      "STORE_total_602_data_0",
      "STORE_total_602_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      STORE_total_573_store_0_req_0,
      STORE_total_573_store_0_ack_0,
      STORE_total_573_store_0_req_1,
      STORE_total_573_store_0_ack_1,
      "STORE_total_573_store_0",
      "memory_space_7" ,
      STORE_total_573_data_0,
      STORE_total_573_word_address_0,
      "STORE_total_573_data_0",
      "STORE_total_573_word_address_0" -- 
    );
    -- shared store operator group (1) : STORE_total_602_store_0 STORE_total_573_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(1 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 7, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 4);
      -- 
    begin -- 
      reqL_unguarded(1) <= STORE_total_602_store_0_req_0;
      reqL_unguarded(0) <= STORE_total_573_store_0_req_0;
      STORE_total_602_store_0_ack_0 <= ackL_unguarded(1);
      STORE_total_573_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= STORE_total_602_store_0_req_1;
      reqR_unguarded(0) <= STORE_total_573_store_0_req_1;
      STORE_total_602_store_0_ack_1 <= ackR_unguarded(1);
      STORE_total_573_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_total_602_word_address_0 & STORE_total_573_word_address_0;
      data_in <= STORE_total_602_data_0 & STORE_total_573_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_7_sr_req(0),
          mack => memory_space_7_sr_ack(0),
          maddr => memory_space_7_sr_addr(0 downto 0),
          mdata => memory_space_7_sr_data(15 downto 0),
          mtag => memory_space_7_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_7_sc_req(0),
          mack => memory_space_7_sc_ack(0),
          mtag => memory_space_7_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- logger for split-operator array_obj_ref_391_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_391_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_391_store_0:started:   inputs: " & " array_obj_ref_391_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_391_word_address_0) & " array_obj_ref_391_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_391_data_0));
          --
        end if; 
        if array_obj_ref_391_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_391_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_398_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_398_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_398_store_0:started:   inputs: " & " array_obj_ref_398_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_398_word_address_0) & " array_obj_ref_398_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_398_data_0));
          --
        end if; 
        if array_obj_ref_398_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_398_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_423_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_423_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_423_store_0:started:   inputs: " & " array_obj_ref_423_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_423_word_address_0) & " array_obj_ref_423_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_423_data_0));
          --
        end if; 
        if array_obj_ref_423_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_423_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_430_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_430_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_430_store_0:started:   inputs: " & " array_obj_ref_430_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_430_word_address_0) & " array_obj_ref_430_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_430_data_0));
          --
        end if; 
        if array_obj_ref_430_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_430_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_391_store_0_req_0,
      array_obj_ref_391_store_0_ack_0,
      array_obj_ref_391_store_0_req_1,
      array_obj_ref_391_store_0_ack_1,
      "array_obj_ref_391_store_0",
      "memory_space_4" ,
      array_obj_ref_391_data_0,
      array_obj_ref_391_word_address_0,
      "array_obj_ref_391_data_0",
      "array_obj_ref_391_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_398_store_0_req_0,
      array_obj_ref_398_store_0_ack_0,
      array_obj_ref_398_store_0_req_1,
      array_obj_ref_398_store_0_ack_1,
      "array_obj_ref_398_store_0",
      "memory_space_4" ,
      array_obj_ref_398_data_0,
      array_obj_ref_398_word_address_0,
      "array_obj_ref_398_data_0",
      "array_obj_ref_398_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_423_store_0_req_0,
      array_obj_ref_423_store_0_ack_0,
      array_obj_ref_423_store_0_req_1,
      array_obj_ref_423_store_0_ack_1,
      "array_obj_ref_423_store_0",
      "memory_space_4" ,
      array_obj_ref_423_data_0,
      array_obj_ref_423_word_address_0,
      "array_obj_ref_423_data_0",
      "array_obj_ref_423_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_430_store_0_req_0,
      array_obj_ref_430_store_0_ack_0,
      array_obj_ref_430_store_0_req_1,
      array_obj_ref_430_store_0_ack_1,
      "array_obj_ref_430_store_0",
      "memory_space_4" ,
      array_obj_ref_430_data_0,
      array_obj_ref_430_word_address_0,
      "array_obj_ref_430_data_0",
      "array_obj_ref_430_word_address_0" -- 
    );
    -- shared store operator group (2) : array_obj_ref_391_store_0 array_obj_ref_398_store_0 array_obj_ref_423_store_0 array_obj_ref_430_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(15 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 7, 2 => 7, 1 => 7, 0 => 7);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 4, 1 => 4, 2 => 4, 3 => 4);
      -- 
    begin -- 
      reqL_unguarded(3) <= array_obj_ref_391_store_0_req_0;
      reqL_unguarded(2) <= array_obj_ref_398_store_0_req_0;
      reqL_unguarded(1) <= array_obj_ref_423_store_0_req_0;
      reqL_unguarded(0) <= array_obj_ref_430_store_0_req_0;
      array_obj_ref_391_store_0_ack_0 <= ackL_unguarded(3);
      array_obj_ref_398_store_0_ack_0 <= ackL_unguarded(2);
      array_obj_ref_423_store_0_ack_0 <= ackL_unguarded(1);
      array_obj_ref_430_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= array_obj_ref_391_store_0_req_1;
      reqR_unguarded(2) <= array_obj_ref_398_store_0_req_1;
      reqR_unguarded(1) <= array_obj_ref_423_store_0_req_1;
      reqR_unguarded(0) <= array_obj_ref_430_store_0_req_1;
      array_obj_ref_391_store_0_ack_1 <= ackR_unguarded(3);
      array_obj_ref_398_store_0_ack_1 <= ackR_unguarded(2);
      array_obj_ref_423_store_0_ack_1 <= ackR_unguarded(1);
      array_obj_ref_430_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      StoreGroup2_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup2_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup2_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_2", num_slots => 2) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup2_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_3", num_slots => 2) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_391_word_address_0 & array_obj_ref_398_word_address_0 & array_obj_ref_423_word_address_0 & array_obj_ref_430_word_address_0;
      data_in <= array_obj_ref_391_data_0 & array_obj_ref_398_data_0 & array_obj_ref_423_data_0 & array_obj_ref_430_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 4,
        data_width => 16,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(3 downto 0),
          mdata => memory_space_4_sr_data(15 downto 0),
          mtag => memory_space_4_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 4,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- logger for split-operator array_obj_ref_547_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_547_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_547_store_0:started:   inputs: " & " array_obj_ref_547_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_547_word_address_0) & " array_obj_ref_547_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_547_data_0));
          --
        end if; 
        if array_obj_ref_547_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_547_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_508_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_508_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_508_store_0:started:   inputs: " & " array_obj_ref_508_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_508_word_address_0) & " array_obj_ref_508_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_508_data_0));
          --
        end if; 
        if array_obj_ref_508_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_508_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_540_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_540_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_540_store_0:started:   inputs: " & " array_obj_ref_540_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_540_word_address_0) & " array_obj_ref_540_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_540_data_0));
          --
        end if; 
        if array_obj_ref_540_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_540_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_657_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_657_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_657_store_0:started:   inputs: " & " array_obj_ref_657_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_657_word_address_0) & " array_obj_ref_657_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_657_data_0));
          --
        end if; 
        if array_obj_ref_657_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_657_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_670_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_670_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_670_store_0:started:   inputs: " & " array_obj_ref_670_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_670_word_address_0) & " array_obj_ref_670_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_670_data_0));
          --
        end if; 
        if array_obj_ref_670_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_670_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_717_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_717_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_717_store_0:started:   inputs: " & " array_obj_ref_717_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_717_word_address_0) & " array_obj_ref_717_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_717_data_0));
          --
        end if; 
        if array_obj_ref_717_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_717_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_683_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_683_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_683_store_0:started:   inputs: " & " array_obj_ref_683_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_683_word_address_0) & " array_obj_ref_683_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_683_data_0));
          --
        end if; 
        if array_obj_ref_683_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_683_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_722_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_722_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_722_store_0:started:   inputs: " & " array_obj_ref_722_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_722_word_address_0) & " array_obj_ref_722_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_722_data_0));
          --
        end if; 
        if array_obj_ref_722_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_722_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_712_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_712_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_712_store_0:started:   inputs: " & " array_obj_ref_712_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_712_word_address_0) & " array_obj_ref_712_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_712_data_0));
          --
        end if; 
        if array_obj_ref_712_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_712_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_707_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_707_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_707_store_0:started:   inputs: " & " array_obj_ref_707_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_707_word_address_0) & " array_obj_ref_707_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_707_data_0));
          --
        end if; 
        if array_obj_ref_707_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_707_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_515_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_515_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_515_store_0:started:   inputs: " & " array_obj_ref_515_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_515_word_address_0) & " array_obj_ref_515_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_515_data_0));
          --
        end if; 
        if array_obj_ref_515_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_515_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_547_store_0_req_0,
      array_obj_ref_547_store_0_ack_0,
      array_obj_ref_547_store_0_req_1,
      array_obj_ref_547_store_0_ack_1,
      "array_obj_ref_547_store_0",
      "memory_space_3" ,
      array_obj_ref_547_data_0,
      array_obj_ref_547_word_address_0,
      "array_obj_ref_547_data_0",
      "array_obj_ref_547_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_508_store_0_req_0,
      array_obj_ref_508_store_0_ack_0,
      array_obj_ref_508_store_0_req_1,
      array_obj_ref_508_store_0_ack_1,
      "array_obj_ref_508_store_0",
      "memory_space_3" ,
      array_obj_ref_508_data_0,
      array_obj_ref_508_word_address_0,
      "array_obj_ref_508_data_0",
      "array_obj_ref_508_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_540_store_0_req_0,
      array_obj_ref_540_store_0_ack_0,
      array_obj_ref_540_store_0_req_1,
      array_obj_ref_540_store_0_ack_1,
      "array_obj_ref_540_store_0",
      "memory_space_3" ,
      array_obj_ref_540_data_0,
      array_obj_ref_540_word_address_0,
      "array_obj_ref_540_data_0",
      "array_obj_ref_540_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_657_store_0_req_0,
      array_obj_ref_657_store_0_ack_0,
      array_obj_ref_657_store_0_req_1,
      array_obj_ref_657_store_0_ack_1,
      "array_obj_ref_657_store_0",
      "memory_space_3" ,
      array_obj_ref_657_data_0,
      array_obj_ref_657_word_address_0,
      "array_obj_ref_657_data_0",
      "array_obj_ref_657_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_670_store_0_req_0,
      array_obj_ref_670_store_0_ack_0,
      array_obj_ref_670_store_0_req_1,
      array_obj_ref_670_store_0_ack_1,
      "array_obj_ref_670_store_0",
      "memory_space_3" ,
      array_obj_ref_670_data_0,
      array_obj_ref_670_word_address_0,
      "array_obj_ref_670_data_0",
      "array_obj_ref_670_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_717_store_0_req_0,
      array_obj_ref_717_store_0_ack_0,
      array_obj_ref_717_store_0_req_1,
      array_obj_ref_717_store_0_ack_1,
      "array_obj_ref_717_store_0",
      "memory_space_3" ,
      array_obj_ref_717_data_0,
      array_obj_ref_717_word_address_0,
      "array_obj_ref_717_data_0",
      "array_obj_ref_717_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_683_store_0_req_0,
      array_obj_ref_683_store_0_ack_0,
      array_obj_ref_683_store_0_req_1,
      array_obj_ref_683_store_0_ack_1,
      "array_obj_ref_683_store_0",
      "memory_space_3" ,
      array_obj_ref_683_data_0,
      array_obj_ref_683_word_address_0,
      "array_obj_ref_683_data_0",
      "array_obj_ref_683_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_722_store_0_req_0,
      array_obj_ref_722_store_0_ack_0,
      array_obj_ref_722_store_0_req_1,
      array_obj_ref_722_store_0_ack_1,
      "array_obj_ref_722_store_0",
      "memory_space_3" ,
      array_obj_ref_722_data_0,
      array_obj_ref_722_word_address_0,
      "array_obj_ref_722_data_0",
      "array_obj_ref_722_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_712_store_0_req_0,
      array_obj_ref_712_store_0_ack_0,
      array_obj_ref_712_store_0_req_1,
      array_obj_ref_712_store_0_ack_1,
      "array_obj_ref_712_store_0",
      "memory_space_3" ,
      array_obj_ref_712_data_0,
      array_obj_ref_712_word_address_0,
      "array_obj_ref_712_data_0",
      "array_obj_ref_712_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_707_store_0_req_0,
      array_obj_ref_707_store_0_ack_0,
      array_obj_ref_707_store_0_req_1,
      array_obj_ref_707_store_0_ack_1,
      "array_obj_ref_707_store_0",
      "memory_space_3" ,
      array_obj_ref_707_data_0,
      array_obj_ref_707_word_address_0,
      "array_obj_ref_707_data_0",
      "array_obj_ref_707_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_515_store_0_req_0,
      array_obj_ref_515_store_0_ack_0,
      array_obj_ref_515_store_0_req_1,
      array_obj_ref_515_store_0_ack_1,
      "array_obj_ref_515_store_0",
      "memory_space_3" ,
      array_obj_ref_515_data_0,
      array_obj_ref_515_word_address_0,
      "array_obj_ref_515_data_0",
      "array_obj_ref_515_word_address_0" -- 
    );
    -- shared store operator group (3) : array_obj_ref_547_store_0 array_obj_ref_508_store_0 array_obj_ref_540_store_0 array_obj_ref_657_store_0 array_obj_ref_670_store_0 array_obj_ref_717_store_0 array_obj_ref_683_store_0 array_obj_ref_722_store_0 array_obj_ref_712_store_0 array_obj_ref_707_store_0 array_obj_ref_515_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(43 downto 0);
      signal data_in: std_logic_vector(175 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 10 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 10 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 10 downto 0);
      signal guard_vector : std_logic_vector( 10 downto 0);
      constant inBUFs : IntegerArray(10 downto 0) := (10 => 2, 9 => 2, 8 => 2, 7 => 2, 6 => 2, 5 => 0, 4 => 2, 3 => 0, 2 => 0, 1 => 0, 0 => 2);
      constant outBUFs : IntegerArray(10 downto 0) := (10 => 7, 9 => 7, 8 => 7, 7 => 7, 6 => 7, 5 => 1, 4 => 7, 3 => 1, 2 => 1, 1 => 1, 0 => 7);
      constant guardFlags : BooleanArray(10 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false);
      constant guardBuffering: IntegerArray(10 downto 0)  := (0 => 4, 1 => 2, 2 => 2, 3 => 2, 4 => 4, 5 => 2, 6 => 4, 7 => 4, 8 => 4, 9 => 4, 10 => 4);
      -- 
    begin -- 
      reqL_unguarded(10) <= array_obj_ref_547_store_0_req_0;
      reqL_unguarded(9) <= array_obj_ref_508_store_0_req_0;
      reqL_unguarded(8) <= array_obj_ref_540_store_0_req_0;
      reqL_unguarded(7) <= array_obj_ref_657_store_0_req_0;
      reqL_unguarded(6) <= array_obj_ref_670_store_0_req_0;
      reqL_unguarded(5) <= array_obj_ref_717_store_0_req_0;
      reqL_unguarded(4) <= array_obj_ref_683_store_0_req_0;
      reqL_unguarded(3) <= array_obj_ref_722_store_0_req_0;
      reqL_unguarded(2) <= array_obj_ref_712_store_0_req_0;
      reqL_unguarded(1) <= array_obj_ref_707_store_0_req_0;
      reqL_unguarded(0) <= array_obj_ref_515_store_0_req_0;
      array_obj_ref_547_store_0_ack_0 <= ackL_unguarded(10);
      array_obj_ref_508_store_0_ack_0 <= ackL_unguarded(9);
      array_obj_ref_540_store_0_ack_0 <= ackL_unguarded(8);
      array_obj_ref_657_store_0_ack_0 <= ackL_unguarded(7);
      array_obj_ref_670_store_0_ack_0 <= ackL_unguarded(6);
      array_obj_ref_717_store_0_ack_0 <= ackL_unguarded(5);
      array_obj_ref_683_store_0_ack_0 <= ackL_unguarded(4);
      array_obj_ref_722_store_0_ack_0 <= ackL_unguarded(3);
      array_obj_ref_712_store_0_ack_0 <= ackL_unguarded(2);
      array_obj_ref_707_store_0_ack_0 <= ackL_unguarded(1);
      array_obj_ref_515_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(10) <= array_obj_ref_547_store_0_req_1;
      reqR_unguarded(9) <= array_obj_ref_508_store_0_req_1;
      reqR_unguarded(8) <= array_obj_ref_540_store_0_req_1;
      reqR_unguarded(7) <= array_obj_ref_657_store_0_req_1;
      reqR_unguarded(6) <= array_obj_ref_670_store_0_req_1;
      reqR_unguarded(5) <= array_obj_ref_717_store_0_req_1;
      reqR_unguarded(4) <= array_obj_ref_683_store_0_req_1;
      reqR_unguarded(3) <= array_obj_ref_722_store_0_req_1;
      reqR_unguarded(2) <= array_obj_ref_712_store_0_req_1;
      reqR_unguarded(1) <= array_obj_ref_707_store_0_req_1;
      reqR_unguarded(0) <= array_obj_ref_515_store_0_req_1;
      array_obj_ref_547_store_0_ack_1 <= ackR_unguarded(10);
      array_obj_ref_508_store_0_ack_1 <= ackR_unguarded(9);
      array_obj_ref_540_store_0_ack_1 <= ackR_unguarded(8);
      array_obj_ref_657_store_0_ack_1 <= ackR_unguarded(7);
      array_obj_ref_670_store_0_ack_1 <= ackR_unguarded(6);
      array_obj_ref_717_store_0_ack_1 <= ackR_unguarded(5);
      array_obj_ref_683_store_0_ack_1 <= ackR_unguarded(4);
      array_obj_ref_722_store_0_ack_1 <= ackR_unguarded(3);
      array_obj_ref_712_store_0_ack_1 <= ackR_unguarded(2);
      array_obj_ref_707_store_0_ack_1 <= ackR_unguarded(1);
      array_obj_ref_515_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      StoreGroup3_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_4: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_4", num_slots => 2) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_5: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_6: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_6", num_slots => 2) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_7: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_7", num_slots => 2) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_8: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_8", num_slots => 2) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_9: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_9", num_slots => 2) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_10: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_10", num_slots => 2) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      StoreGroup3_gI: SplitGuardInterface generic map(name => "StoreGroup3_gI", nreqs => 11, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_547_word_address_0 & array_obj_ref_508_word_address_0 & array_obj_ref_540_word_address_0 & array_obj_ref_657_word_address_0 & array_obj_ref_670_word_address_0 & array_obj_ref_717_word_address_0 & array_obj_ref_683_word_address_0 & array_obj_ref_722_word_address_0 & array_obj_ref_712_word_address_0 & array_obj_ref_707_word_address_0 & array_obj_ref_515_word_address_0;
      data_in <= array_obj_ref_547_data_0 & array_obj_ref_508_data_0 & array_obj_ref_540_data_0 & array_obj_ref_657_data_0 & array_obj_ref_670_data_0 & array_obj_ref_717_data_0 & array_obj_ref_683_data_0 & array_obj_ref_722_data_0 & array_obj_ref_712_data_0 & array_obj_ref_707_data_0 & array_obj_ref_515_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup3 Req ", addr_width => 4,
        data_width => 16,
        num_reqs => 11,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(3 downto 0),
          mdata => memory_space_3_sr_data(15 downto 0),
          mtag => memory_space_3_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup3 Complete ",
          num_reqs => 11,
          detailed_buffering_per_output => outBUFs,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- logger for split-operator array_obj_ref_597_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_597_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_597_store_0:started:   inputs: " & " array_obj_ref_597_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_597_word_address_0) & " array_obj_ref_597_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_597_data_0));
          --
        end if; 
        if array_obj_ref_597_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:array_obj_ref_597_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_597_store_0_req_0,
      array_obj_ref_597_store_0_ack_0,
      array_obj_ref_597_store_0_req_1,
      array_obj_ref_597_store_0_ack_1,
      "array_obj_ref_597_store_0",
      "memory_space_2" ,
      array_obj_ref_597_data_0,
      array_obj_ref_597_word_address_0,
      "array_obj_ref_597_data_0",
      "array_obj_ref_597_word_address_0" -- 
    );
    -- shared store operator group (4) : array_obj_ref_597_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(3 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 7);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_597_store_0_req_0;
      array_obj_ref_597_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_597_store_0_req_1;
      array_obj_ref_597_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup4_gI: SplitGuardInterface generic map(name => "StoreGroup4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_597_word_address_0;
      data_in <= array_obj_ref_597_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup4 Req ", addr_width => 4,
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(3 downto 0),
          mdata => memory_space_2_sr_data(15 downto 0),
          mtag => memory_space_2_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup4 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- logger for split-operator WPIPE_acc_mem_635_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_acc_mem_635_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:WPIPE_acc_mem_635_inst:started:   PipeWrite to acc_mem inputs: " & " array_obj_ref_637_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_637_wire));
          --
        end if; 
        if WPIPE_acc_mem_635_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:WPIPE_acc_mem_635_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_acc_mem_635_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_acc_mem_635_inst_req_0;
      WPIPE_acc_mem_635_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_acc_mem_635_inst_req_1;
      WPIPE_acc_mem_635_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= array_obj_ref_637_wire;
      acc_mem_write_0_gI: SplitGuardInterface generic map(name => "acc_mem_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      acc_mem_write_0: OutputPortRevised -- 
        generic map ( name => "acc_mem", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => acc_mem_pipe_write_req(0),
          oack => acc_mem_pipe_write_ack(0),
          odata => acc_mem_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logger for split-operator WPIPE_acc_mem_add_632_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_acc_mem_add_632_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:WPIPE_acc_mem_add_632_inst:started:   PipeWrite to acc_mem_add inputs: " & " f_631 = "& Convert_SLV_To_Hex_String(f_631));
          --
        end if; 
        if WPIPE_acc_mem_add_632_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:WPIPE_acc_mem_add_632_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (1) : WPIPE_acc_mem_add_632_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_acc_mem_add_632_inst_req_0;
      WPIPE_acc_mem_add_632_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_acc_mem_add_632_inst_req_1;
      WPIPE_acc_mem_add_632_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= f_631;
      acc_mem_add_write_1_gI: SplitGuardInterface generic map(name => "acc_mem_add_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      acc_mem_add_write_1: OutputPortRevised -- 
        generic map ( name => "acc_mem_add", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => acc_mem_add_pipe_write_req(0),
          oack => acc_mem_add_pipe_write_ack(0),
          odata => acc_mem_add_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- logger for split-operator call_stmt_373_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_373_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:call_stmt_373_call:started:  Call to module accMemAccessDaemon inputs: " & " NNT_369 = "& Convert_SLV_To_Hex_String(NNT_369));
          --
        end if; 
        if call_stmt_373_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:call_stmt_373_call:finished:  outputs: " & " rdatalk_373= "  & Convert_SLV_To_Hex_String(rdatalk_373) & " rdatahk_373= "  & Convert_SLV_To_Hex_String(rdatahk_373));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_490_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_490_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:call_stmt_490_call:started:  Call to module accMemAccessDaemon inputs: " & " NNJ_486 = "& Convert_SLV_To_Hex_String(NNJ_486));
          --
        end if; 
        if call_stmt_490_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:call_stmt_490_call:finished:  outputs: " & " rdatal_490= "  & Convert_SLV_To_Hex_String(rdatal_490) & " rdatah_490= "  & Convert_SLV_To_Hex_String(rdatah_490));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_373_call call_stmt_490_call 
    accMemAccessDaemon_call_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 4, 1 => 4);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_373_call_req_0;
      reqL_unguarded(0) <= call_stmt_490_call_req_0;
      call_stmt_373_call_ack_0 <= ackL_unguarded(1);
      call_stmt_490_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_373_call_req_1;
      reqR_unguarded(0) <= call_stmt_490_call_req_1;
      call_stmt_373_call_ack_1 <= ackR_unguarded(1);
      call_stmt_490_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accMemAccessDaemon_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accMemAccessDaemon_call_group_0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accMemAccessDaemon_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accMemAccessDaemon_call_group_0_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accMemAccessDaemon_call_group_0_gI: SplitGuardInterface generic map(name => "accMemAccessDaemon_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= NNT_369 & NNJ_486;
      rdatalk_373 <= data_out(127 downto 96);
      rdatahk_373 <= data_out(95 downto 64);
      rdatal_490 <= data_out(63 downto 32);
      rdatah_490 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 64,
        owidth => 32,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accMemAccessDaemon_call_reqs(0),
          ackR => accMemAccessDaemon_call_acks(0),
          dataR => accMemAccessDaemon_call_data(31 downto 0),
          tagR => accMemAccessDaemon_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accMemAccessDaemon_return_acks(0), -- cross-over
          ackL => accMemAccessDaemon_return_reqs(0), -- cross-over
          dataL => accMemAccessDaemon_return_data(63 downto 0),
          tagL => accMemAccessDaemon_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- logger for split-operator call_stmt_624_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_624_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:call_stmt_624_call:started:  Call to module accessMem inputs: " & " konst_618_wire_constant = "& Convert_SLV_To_Hex_String(konst_618_wire_constant) & " ADD_u12_u12_621_wire = "& Convert_SLV_To_Hex_String(ADD_u12_u12_621_wire) & " LOAD_total_622_wire = "& Convert_SLV_To_Hex_String(LOAD_total_622_wire));
          --
        end if; 
        if call_stmt_624_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:call_stmt_624_call:finished:  outputs: " & " rdata_624= "  & Convert_SLV_To_Hex_String(rdata_624));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (1) : call_stmt_624_call 
    accessMem_call_group_1: Block -- 
      signal data_in: std_logic_vector(28 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_624_call_req_0;
      call_stmt_624_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_624_call_req_1;
      call_stmt_624_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMem_call_group_1_gI: SplitGuardInterface generic map(name => "accessMem_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_618_wire_constant & ADD_u12_u12_621_wire & LOAD_total_622_wire;
      rdata_624 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 29,
        owidth => 29,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMem_call_reqs(0),
          ackR => accessMem_call_acks(0),
          dataR => accessMem_call_data(28 downto 0),
          tagR => accessMem_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMem_return_acks(0), -- cross-over
          ackL => accessMem_return_reqs(0), -- cross-over
          dataL => accessMem_return_data(63 downto 0),
          tagL => accessMem_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- logger for split-operator call_stmt_705_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_705_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:call_stmt_705_call:started:  Call to module accessMem_v inputs: " & " konst_697_wire_constant = "& Convert_SLV_To_Hex_String(konst_697_wire_constant) & " ADD_u12_u12_702_wire = "& Convert_SLV_To_Hex_String(ADD_u12_u12_702_wire) & " konst_703_wire_constant = "& Convert_SLV_To_Hex_String(konst_703_wire_constant));
          --
        end if; 
        if call_stmt_705_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:try1:DP:call_stmt_705_call:finished:  outputs: " & " rdatar_705= "  & Convert_SLV_To_Hex_String(rdatar_705));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (2) : call_stmt_705_call 
    accessMem_v_call_group_2: Block -- 
      signal data_in: std_logic_vector(28 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_705_call_req_0;
      call_stmt_705_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_705_call_req_1;
      call_stmt_705_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMem_v_call_group_2_gI: SplitGuardInterface generic map(name => "accessMem_v_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_697_wire_constant & ADD_u12_u12_702_wire & konst_703_wire_constant;
      rdatar_705 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 29,
        owidth => 29,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMem_v_call_reqs(0),
          ackR => accessMem_v_call_acks(0),
          dataR => accessMem_v_call_data(28 downto 0),
          tagR => accessMem_v_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMem_v_return_acks(0), -- cross-over
          ackL => accessMem_v_return_reqs(0), -- cross-over
          dataL => accessMem_v_return_data(63 downto 0),
          tagL => accessMem_v_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end try1_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    acc_mem_pipe_read_data: out std_logic_vector(15 downto 0);
    acc_mem_pipe_read_req : in std_logic_vector(0 downto 0);
    acc_mem_pipe_read_ack : out std_logic_vector(0 downto 0);
    acc_mem_add_pipe_read_data: out std_logic_vector(15 downto 0);
    acc_mem_add_pipe_read_req : in std_logic_vector(0 downto 0);
    acc_mem_add_pipe_read_ack : out std_logic_vector(0 downto 0);
    start_pipe_write_data: in std_logic_vector(15 downto 0);
    start_pipe_write_req : in std_logic_vector(0 downto 0);
    start_pipe_write_ack : out std_logic_vector(0 downto 0);
    status_pipe_read_data: out std_logic_vector(15 downto 0);
    status_pipe_read_req : in std_logic_vector(0 downto 0);
    status_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(1 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(37 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(23 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(11 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(3 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(3 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(20 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_lr_addr : std_logic_vector(3 downto 0);
  signal memory_space_4_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_4_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_4_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_4_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_5
  signal memory_space_5_lr_req :  std_logic_vector(2 downto 0);
  signal memory_space_5_lr_ack : std_logic_vector(2 downto 0);
  signal memory_space_5_lr_addr : std_logic_vector(32 downto 0);
  signal memory_space_5_lr_tag : std_logic_vector(62 downto 0);
  signal memory_space_5_lc_req : std_logic_vector(2 downto 0);
  signal memory_space_5_lc_ack :  std_logic_vector(2 downto 0);
  signal memory_space_5_lc_data : std_logic_vector(47 downto 0);
  signal memory_space_5_lc_tag :  std_logic_vector(8 downto 0);
  signal memory_space_5_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_5_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_5_sr_addr : std_logic_vector(21 downto 0);
  signal memory_space_5_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_5_sr_tag : std_logic_vector(41 downto 0);
  signal memory_space_5_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_5_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_5_sc_tag :  std_logic_vector(5 downto 0);
  -- interface signals to connect to memory space memory_space_6
  signal memory_space_6_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_6_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_6_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_lc_data : std_logic_vector(0 downto 0);
  signal memory_space_6_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_6_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_data : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_6_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_7
  signal memory_space_7_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_7_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_7_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_7_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_7_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_7_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_8
  signal memory_space_8_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_8_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_8_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_8_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_8_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_8_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_8_lc_data : std_logic_vector(3 downto 0);
  signal memory_space_8_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_8_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_8_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_data : std_logic_vector(3 downto 0);
  signal memory_space_8_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_8_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_8_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_8_sc_tag :  std_logic_vector(0 downto 0);
  -- declarations related to module accMemAccessDaemon
  component accMemAccessDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      acc_mem_request : in  std_logic_vector(31 downto 0);
      acc_mem_responsel : out  std_logic_vector(31 downto 0);
      acc_mem_responseh : out  std_logic_vector(31 downto 0);
      accessMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessMem_call_acks : in   std_logic_vector(0 downto 0);
      accessMem_call_data : out  std_logic_vector(28 downto 0);
      accessMem_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessMem_return_acks : in   std_logic_vector(0 downto 0);
      accessMem_return_data : in   std_logic_vector(63 downto 0);
      accessMem_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accMemAccessDaemon
  signal accMemAccessDaemon_acc_mem_request :  std_logic_vector(31 downto 0);
  signal accMemAccessDaemon_acc_mem_responsel :  std_logic_vector(31 downto 0);
  signal accMemAccessDaemon_acc_mem_responseh :  std_logic_vector(31 downto 0);
  signal accMemAccessDaemon_in_args    : std_logic_vector(31 downto 0);
  signal accMemAccessDaemon_out_args   : std_logic_vector(63 downto 0);
  signal accMemAccessDaemon_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal accMemAccessDaemon_tag_out   : std_logic_vector(2 downto 0);
  signal accMemAccessDaemon_start_req : std_logic;
  signal accMemAccessDaemon_start_ack : std_logic;
  signal accMemAccessDaemon_fin_req   : std_logic;
  signal accMemAccessDaemon_fin_ack : std_logic;
  -- caller side aggregated signals for module accMemAccessDaemon
  signal accMemAccessDaemon_call_reqs: std_logic_vector(0 downto 0);
  signal accMemAccessDaemon_call_acks: std_logic_vector(0 downto 0);
  signal accMemAccessDaemon_return_reqs: std_logic_vector(0 downto 0);
  signal accMemAccessDaemon_return_acks: std_logic_vector(0 downto 0);
  signal accMemAccessDaemon_call_data: std_logic_vector(31 downto 0);
  signal accMemAccessDaemon_call_tag: std_logic_vector(1 downto 0);
  signal accMemAccessDaemon_return_data: std_logic_vector(63 downto 0);
  signal accMemAccessDaemon_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module accessMem
  component accessMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(11 downto 0);
      write_data : in  std_logic_vector(15 downto 0);
      read_datal : out  std_logic_vector(63 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessMem
  signal accessMem_read_write_bar :  std_logic_vector(0 downto 0);
  signal accessMem_addr :  std_logic_vector(11 downto 0);
  signal accessMem_write_data :  std_logic_vector(15 downto 0);
  signal accessMem_read_datal :  std_logic_vector(63 downto 0);
  signal accessMem_in_args    : std_logic_vector(28 downto 0);
  signal accessMem_out_args   : std_logic_vector(63 downto 0);
  signal accessMem_tag_in    : std_logic_vector(4 downto 0) := (others => '0');
  signal accessMem_tag_out   : std_logic_vector(4 downto 0);
  signal accessMem_start_req : std_logic;
  signal accessMem_start_ack : std_logic;
  signal accessMem_fin_req   : std_logic;
  signal accessMem_fin_ack : std_logic;
  -- caller side aggregated signals for module accessMem
  signal accessMem_call_reqs: std_logic_vector(4 downto 0);
  signal accessMem_call_acks: std_logic_vector(4 downto 0);
  signal accessMem_return_reqs: std_logic_vector(4 downto 0);
  signal accessMem_return_acks: std_logic_vector(4 downto 0);
  signal accessMem_call_data: std_logic_vector(144 downto 0);
  signal accessMem_call_tag: std_logic_vector(9 downto 0);
  signal accessMem_return_data: std_logic_vector(319 downto 0);
  signal accessMem_return_tag: std_logic_vector(9 downto 0);
  -- declarations related to module accessMem_v
  component accessMem_v is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(11 downto 0);
      write_data : in  std_logic_vector(15 downto 0);
      read_datal : out  std_logic_vector(63 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessMem_v
  signal accessMem_v_read_write_bar :  std_logic_vector(0 downto 0);
  signal accessMem_v_addr :  std_logic_vector(11 downto 0);
  signal accessMem_v_write_data :  std_logic_vector(15 downto 0);
  signal accessMem_v_read_datal :  std_logic_vector(63 downto 0);
  signal accessMem_v_in_args    : std_logic_vector(28 downto 0);
  signal accessMem_v_out_args   : std_logic_vector(63 downto 0);
  signal accessMem_v_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal accessMem_v_tag_out   : std_logic_vector(1 downto 0);
  signal accessMem_v_start_req : std_logic;
  signal accessMem_v_start_ack : std_logic;
  signal accessMem_v_fin_req   : std_logic;
  signal accessMem_v_fin_ack : std_logic;
  -- caller side aggregated signals for module accessMem_v
  signal accessMem_v_call_reqs: std_logic_vector(0 downto 0);
  signal accessMem_v_call_acks: std_logic_vector(0 downto 0);
  signal accessMem_v_return_reqs: std_logic_vector(0 downto 0);
  signal accessMem_v_return_acks: std_logic_vector(0 downto 0);
  signal accessMem_v_call_data: std_logic_vector(28 downto 0);
  signal accessMem_v_call_tag: std_logic_vector(0 downto 0);
  signal accessMem_v_return_data: std_logic_vector(63 downto 0);
  signal accessMem_v_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module initial
  component initial is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(11 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(11 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      accessMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessMem_call_acks : in   std_logic_vector(0 downto 0);
      accessMem_call_data : out  std_logic_vector(28 downto 0);
      accessMem_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessMem_return_acks : in   std_logic_vector(0 downto 0);
      accessMem_return_data : in   std_logic_vector(63 downto 0);
      accessMem_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module initial
  signal initial_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal initial_tag_out   : std_logic_vector(1 downto 0);
  signal initial_start_req : std_logic;
  signal initial_start_ack : std_logic;
  signal initial_fin_req   : std_logic;
  signal initial_fin_ack : std_logic;
  -- caller side aggregated signals for module initial
  signal initial_call_reqs: std_logic_vector(0 downto 0);
  signal initial_call_acks: std_logic_vector(0 downto 0);
  signal initial_return_reqs: std_logic_vector(0 downto 0);
  signal initial_return_acks: std_logic_vector(0 downto 0);
  signal initial_call_tag: std_logic_vector(0 downto 0);
  signal initial_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module try
  component try is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(3 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(0 downto 0);
      start_pipe_read_req : out  std_logic_vector(0 downto 0);
      start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      start_pipe_read_data : in   std_logic_vector(15 downto 0);
      status_pipe_write_req : out  std_logic_vector(0 downto 0);
      status_pipe_write_ack : in   std_logic_vector(0 downto 0);
      status_pipe_write_data : out  std_logic_vector(15 downto 0);
      accessMem_call_reqs : out  std_logic_vector(1 downto 0);
      accessMem_call_acks : in   std_logic_vector(1 downto 0);
      accessMem_call_data : out  std_logic_vector(57 downto 0);
      accessMem_call_tag  :  out  std_logic_vector(3 downto 0);
      accessMem_return_reqs : out  std_logic_vector(1 downto 0);
      accessMem_return_acks : in   std_logic_vector(1 downto 0);
      accessMem_return_data : in   std_logic_vector(127 downto 0);
      accessMem_return_tag :  in   std_logic_vector(3 downto 0);
      initial_call_reqs : out  std_logic_vector(0 downto 0);
      initial_call_acks : in   std_logic_vector(0 downto 0);
      initial_call_tag  :  out  std_logic_vector(0 downto 0);
      initial_return_reqs : out  std_logic_vector(0 downto 0);
      initial_return_acks : in   std_logic_vector(0 downto 0);
      initial_return_tag :  in   std_logic_vector(0 downto 0);
      try1_call_reqs : out  std_logic_vector(0 downto 0);
      try1_call_acks : in   std_logic_vector(0 downto 0);
      try1_call_tag  :  out  std_logic_vector(0 downto 0);
      try1_return_reqs : out  std_logic_vector(0 downto 0);
      try1_return_acks : in   std_logic_vector(0 downto 0);
      try1_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module try
  signal try_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal try_tag_out   : std_logic_vector(1 downto 0);
  signal try_start_req : std_logic;
  signal try_start_ack : std_logic;
  signal try_fin_req   : std_logic;
  signal try_fin_ack : std_logic;
  -- declarations related to module try1
  component try1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(11 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(3 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(1 downto 0);
      acc_mem_pipe_write_req : out  std_logic_vector(0 downto 0);
      acc_mem_pipe_write_ack : in   std_logic_vector(0 downto 0);
      acc_mem_pipe_write_data : out  std_logic_vector(15 downto 0);
      acc_mem_add_pipe_write_req : out  std_logic_vector(0 downto 0);
      acc_mem_add_pipe_write_ack : in   std_logic_vector(0 downto 0);
      acc_mem_add_pipe_write_data : out  std_logic_vector(15 downto 0);
      accessMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessMem_call_acks : in   std_logic_vector(0 downto 0);
      accessMem_call_data : out  std_logic_vector(28 downto 0);
      accessMem_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessMem_return_acks : in   std_logic_vector(0 downto 0);
      accessMem_return_data : in   std_logic_vector(63 downto 0);
      accessMem_return_tag :  in   std_logic_vector(1 downto 0);
      accessMem_v_call_reqs : out  std_logic_vector(0 downto 0);
      accessMem_v_call_acks : in   std_logic_vector(0 downto 0);
      accessMem_v_call_data : out  std_logic_vector(28 downto 0);
      accessMem_v_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMem_v_return_reqs : out  std_logic_vector(0 downto 0);
      accessMem_v_return_acks : in   std_logic_vector(0 downto 0);
      accessMem_v_return_data : in   std_logic_vector(63 downto 0);
      accessMem_v_return_tag :  in   std_logic_vector(0 downto 0);
      accMemAccessDaemon_call_reqs : out  std_logic_vector(0 downto 0);
      accMemAccessDaemon_call_acks : in   std_logic_vector(0 downto 0);
      accMemAccessDaemon_call_data : out  std_logic_vector(31 downto 0);
      accMemAccessDaemon_call_tag  :  out  std_logic_vector(1 downto 0);
      accMemAccessDaemon_return_reqs : out  std_logic_vector(0 downto 0);
      accMemAccessDaemon_return_acks : in   std_logic_vector(0 downto 0);
      accMemAccessDaemon_return_data : in   std_logic_vector(63 downto 0);
      accMemAccessDaemon_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module try1
  signal try1_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal try1_tag_out   : std_logic_vector(1 downto 0);
  signal try1_start_req : std_logic;
  signal try1_start_ack : std_logic;
  signal try1_fin_req   : std_logic;
  signal try1_fin_ack : std_logic;
  -- caller side aggregated signals for module try1
  signal try1_call_reqs: std_logic_vector(0 downto 0);
  signal try1_call_acks: std_logic_vector(0 downto 0);
  signal try1_return_reqs: std_logic_vector(0 downto 0);
  signal try1_return_acks: std_logic_vector(0 downto 0);
  signal try1_call_tag: std_logic_vector(0 downto 0);
  signal try1_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe acc_mem
  signal acc_mem_pipe_write_data: std_logic_vector(15 downto 0);
  signal acc_mem_pipe_write_req: std_logic_vector(0 downto 0);
  signal acc_mem_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe acc_mem_add
  signal acc_mem_add_pipe_write_data: std_logic_vector(15 downto 0);
  signal acc_mem_add_pipe_write_req: std_logic_vector(0 downto 0);
  signal acc_mem_add_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe start
  signal start_pipe_read_data: std_logic_vector(15 downto 0);
  signal start_pipe_read_req: std_logic_vector(0 downto 0);
  signal start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe status
  signal status_pipe_write_data: std_logic_vector(15 downto 0);
  signal status_pipe_write_req: std_logic_vector(0 downto 0);
  signal status_pipe_write_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module accMemAccessDaemon
  accMemAccessDaemon_acc_mem_request <= accMemAccessDaemon_in_args(31 downto 0);
  accMemAccessDaemon_out_args <= accMemAccessDaemon_acc_mem_responsel & accMemAccessDaemon_acc_mem_responseh ;
  -- call arbiter for module accMemAccessDaemon
  accMemAccessDaemon_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 32,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => accMemAccessDaemon_call_reqs,
      call_acks => accMemAccessDaemon_call_acks,
      return_reqs => accMemAccessDaemon_return_reqs,
      return_acks => accMemAccessDaemon_return_acks,
      call_data  => accMemAccessDaemon_call_data,
      call_tag  => accMemAccessDaemon_call_tag,
      return_tag  => accMemAccessDaemon_return_tag,
      call_mtag => accMemAccessDaemon_tag_in,
      return_mtag => accMemAccessDaemon_tag_out,
      return_data =>accMemAccessDaemon_return_data,
      call_mreq => accMemAccessDaemon_start_req,
      call_mack => accMemAccessDaemon_start_ack,
      return_mreq => accMemAccessDaemon_fin_req,
      return_mack => accMemAccessDaemon_fin_ack,
      call_mdata => accMemAccessDaemon_in_args,
      return_mdata => accMemAccessDaemon_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accMemAccessDaemon_instance:accMemAccessDaemon-- 
    generic map(tag_length => 3)
    port map(-- 
      acc_mem_request => accMemAccessDaemon_acc_mem_request,
      acc_mem_responsel => accMemAccessDaemon_acc_mem_responsel,
      acc_mem_responseh => accMemAccessDaemon_acc_mem_responseh,
      start_req => accMemAccessDaemon_start_req,
      start_ack => accMemAccessDaemon_start_ack,
      fin_req => accMemAccessDaemon_fin_req,
      fin_ack => accMemAccessDaemon_fin_ack,
      clk => clk,
      reset => reset,
      accessMem_call_reqs => accessMem_call_reqs(3 downto 3),
      accessMem_call_acks => accessMem_call_acks(3 downto 3),
      accessMem_call_data => accessMem_call_data(115 downto 87),
      accessMem_call_tag => accessMem_call_tag(7 downto 6),
      accessMem_return_reqs => accessMem_return_reqs(3 downto 3),
      accessMem_return_acks => accessMem_return_acks(3 downto 3),
      accessMem_return_data => accessMem_return_data(255 downto 192),
      accessMem_return_tag => accessMem_return_tag(7 downto 6),
      tag_in => accMemAccessDaemon_tag_in,
      tag_out => accMemAccessDaemon_tag_out-- 
    ); -- 
  -- module accessMem
  accessMem_read_write_bar <= accessMem_in_args(28 downto 28);
  accessMem_addr <= accessMem_in_args(27 downto 16);
  accessMem_write_data <= accessMem_in_args(15 downto 0);
  accessMem_out_args <= accessMem_read_datal ;
  -- call arbiter for module accessMem
  accessMem_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 5,
      call_data_width => 29,
      return_data_width => 64,
      callee_tag_length => 3,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => accessMem_call_reqs,
      call_acks => accessMem_call_acks,
      return_reqs => accessMem_return_reqs,
      return_acks => accessMem_return_acks,
      call_data  => accessMem_call_data,
      call_tag  => accessMem_call_tag,
      return_tag  => accessMem_return_tag,
      call_mtag => accessMem_tag_in,
      return_mtag => accessMem_tag_out,
      return_data =>accessMem_return_data,
      call_mreq => accessMem_start_req,
      call_mack => accessMem_start_ack,
      return_mreq => accessMem_fin_req,
      return_mack => accessMem_fin_ack,
      call_mdata => accessMem_in_args,
      return_mdata => accessMem_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessMem_instance:accessMem-- 
    generic map(tag_length => 5)
    port map(-- 
      read_write_bar => accessMem_read_write_bar,
      addr => accessMem_addr,
      write_data => accessMem_write_data,
      read_datal => accessMem_read_datal,
      start_req => accessMem_start_req,
      start_ack => accessMem_start_ack,
      fin_req => accessMem_fin_req,
      fin_ack => accessMem_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_lr_req => memory_space_5_lr_req(2 downto 2),
      memory_space_5_lr_ack => memory_space_5_lr_ack(2 downto 2),
      memory_space_5_lr_addr => memory_space_5_lr_addr(32 downto 22),
      memory_space_5_lr_tag => memory_space_5_lr_tag(62 downto 42),
      memory_space_5_lc_req => memory_space_5_lc_req(2 downto 2),
      memory_space_5_lc_ack => memory_space_5_lc_ack(2 downto 2),
      memory_space_5_lc_data => memory_space_5_lc_data(47 downto 32),
      memory_space_5_lc_tag => memory_space_5_lc_tag(8 downto 6),
      memory_space_5_sr_req => memory_space_5_sr_req(1 downto 1),
      memory_space_5_sr_ack => memory_space_5_sr_ack(1 downto 1),
      memory_space_5_sr_addr => memory_space_5_sr_addr(21 downto 11),
      memory_space_5_sr_data => memory_space_5_sr_data(31 downto 16),
      memory_space_5_sr_tag => memory_space_5_sr_tag(41 downto 21),
      memory_space_5_sc_req => memory_space_5_sc_req(1 downto 1),
      memory_space_5_sc_ack => memory_space_5_sc_ack(1 downto 1),
      memory_space_5_sc_tag => memory_space_5_sc_tag(5 downto 3),
      tag_in => accessMem_tag_in,
      tag_out => accessMem_tag_out-- 
    ); -- 
  -- module accessMem_v
  accessMem_v_read_write_bar <= accessMem_v_in_args(28 downto 28);
  accessMem_v_addr <= accessMem_v_in_args(27 downto 16);
  accessMem_v_write_data <= accessMem_v_in_args(15 downto 0);
  accessMem_v_out_args <= accessMem_v_read_datal ;
  -- call arbiter for module accessMem_v
  accessMem_v_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 29,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => accessMem_v_call_reqs,
      call_acks => accessMem_v_call_acks,
      return_reqs => accessMem_v_return_reqs,
      return_acks => accessMem_v_return_acks,
      call_data  => accessMem_v_call_data,
      call_tag  => accessMem_v_call_tag,
      return_tag  => accessMem_v_return_tag,
      call_mtag => accessMem_v_tag_in,
      return_mtag => accessMem_v_tag_out,
      return_data =>accessMem_v_return_data,
      call_mreq => accessMem_v_start_req,
      call_mack => accessMem_v_start_ack,
      return_mreq => accessMem_v_fin_req,
      return_mack => accessMem_v_fin_ack,
      call_mdata => accessMem_v_in_args,
      return_mdata => accessMem_v_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessMem_v_instance:accessMem_v-- 
    generic map(tag_length => 2)
    port map(-- 
      read_write_bar => accessMem_v_read_write_bar,
      addr => accessMem_v_addr,
      write_data => accessMem_v_write_data,
      read_datal => accessMem_v_read_datal,
      start_req => accessMem_v_start_req,
      start_ack => accessMem_v_start_ack,
      fin_req => accessMem_v_fin_req,
      fin_ack => accessMem_v_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_lr_req => memory_space_5_lr_req(1 downto 1),
      memory_space_5_lr_ack => memory_space_5_lr_ack(1 downto 1),
      memory_space_5_lr_addr => memory_space_5_lr_addr(21 downto 11),
      memory_space_5_lr_tag => memory_space_5_lr_tag(41 downto 21),
      memory_space_5_lc_req => memory_space_5_lc_req(1 downto 1),
      memory_space_5_lc_ack => memory_space_5_lc_ack(1 downto 1),
      memory_space_5_lc_data => memory_space_5_lc_data(31 downto 16),
      memory_space_5_lc_tag => memory_space_5_lc_tag(5 downto 3),
      memory_space_5_sr_req => memory_space_5_sr_req(0 downto 0),
      memory_space_5_sr_ack => memory_space_5_sr_ack(0 downto 0),
      memory_space_5_sr_addr => memory_space_5_sr_addr(10 downto 0),
      memory_space_5_sr_data => memory_space_5_sr_data(15 downto 0),
      memory_space_5_sr_tag => memory_space_5_sr_tag(20 downto 0),
      memory_space_5_sc_req => memory_space_5_sc_req(0 downto 0),
      memory_space_5_sc_ack => memory_space_5_sc_ack(0 downto 0),
      memory_space_5_sc_tag => memory_space_5_sc_tag(2 downto 0),
      tag_in => accessMem_v_tag_in,
      tag_out => accessMem_v_tag_out-- 
    ); -- 
  -- module initial
  -- call arbiter for module initial
  initial_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => initial_call_reqs,
      call_acks => initial_call_acks,
      return_reqs => initial_return_reqs,
      return_acks => initial_return_acks,
      call_tag  => initial_call_tag,
      return_tag  => initial_return_tag,
      call_mtag => initial_tag_in,
      return_mtag => initial_tag_out,
      call_mreq => initial_start_req,
      call_mack => initial_start_ack,
      return_mreq => initial_fin_req,
      return_mack => initial_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  initial_instance:initial-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => initial_start_req,
      start_ack => initial_start_ack,
      fin_req => initial_fin_req,
      fin_ack => initial_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(1 downto 1),
      memory_space_1_lr_tag => memory_space_1_lr_tag(37 downto 19),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(23 downto 12),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 2),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(0 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(11 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(1 downto 0),
      accessMem_call_reqs => accessMem_call_reqs(4 downto 4),
      accessMem_call_acks => accessMem_call_acks(4 downto 4),
      accessMem_call_data => accessMem_call_data(144 downto 116),
      accessMem_call_tag => accessMem_call_tag(9 downto 8),
      accessMem_return_reqs => accessMem_return_reqs(4 downto 4),
      accessMem_return_acks => accessMem_return_acks(4 downto 4),
      accessMem_return_data => accessMem_return_data(319 downto 256),
      accessMem_return_tag => accessMem_return_tag(9 downto 8),
      tag_in => initial_tag_in,
      tag_out => initial_tag_out-- 
    ); -- 
  -- module try
  try_instance:try-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => try_start_req,
      start_ack => try_start_ack,
      fin_req => try_fin_req,
      fin_ack => try_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_6_sr_req => memory_space_6_sr_req(0 downto 0),
      memory_space_6_sr_ack => memory_space_6_sr_ack(0 downto 0),
      memory_space_6_sr_addr => memory_space_6_sr_addr(0 downto 0),
      memory_space_6_sr_data => memory_space_6_sr_data(0 downto 0),
      memory_space_6_sr_tag => memory_space_6_sr_tag(18 downto 0),
      memory_space_6_sc_req => memory_space_6_sc_req(0 downto 0),
      memory_space_6_sc_ack => memory_space_6_sc_ack(0 downto 0),
      memory_space_6_sc_tag => memory_space_6_sc_tag(1 downto 0),
      memory_space_8_sr_req => memory_space_8_sr_req(0 downto 0),
      memory_space_8_sr_ack => memory_space_8_sr_ack(0 downto 0),
      memory_space_8_sr_addr => memory_space_8_sr_addr(0 downto 0),
      memory_space_8_sr_data => memory_space_8_sr_data(3 downto 0),
      memory_space_8_sr_tag => memory_space_8_sr_tag(17 downto 0),
      memory_space_8_sc_req => memory_space_8_sc_req(0 downto 0),
      memory_space_8_sc_ack => memory_space_8_sc_ack(0 downto 0),
      memory_space_8_sc_tag => memory_space_8_sc_tag(0 downto 0),
      start_pipe_read_req => start_pipe_read_req(0 downto 0),
      start_pipe_read_ack => start_pipe_read_ack(0 downto 0),
      start_pipe_read_data => start_pipe_read_data(15 downto 0),
      status_pipe_write_req => status_pipe_write_req(0 downto 0),
      status_pipe_write_ack => status_pipe_write_ack(0 downto 0),
      status_pipe_write_data => status_pipe_write_data(15 downto 0),
      accessMem_call_reqs => accessMem_call_reqs(1 downto 0),
      accessMem_call_acks => accessMem_call_acks(1 downto 0),
      accessMem_call_data => accessMem_call_data(57 downto 0),
      accessMem_call_tag => accessMem_call_tag(3 downto 0),
      accessMem_return_reqs => accessMem_return_reqs(1 downto 0),
      accessMem_return_acks => accessMem_return_acks(1 downto 0),
      accessMem_return_data => accessMem_return_data(127 downto 0),
      accessMem_return_tag => accessMem_return_tag(3 downto 0),
      initial_call_reqs => initial_call_reqs(0 downto 0),
      initial_call_acks => initial_call_acks(0 downto 0),
      initial_call_tag => initial_call_tag(0 downto 0),
      initial_return_reqs => initial_return_reqs(0 downto 0),
      initial_return_acks => initial_return_acks(0 downto 0),
      initial_return_tag => initial_return_tag(0 downto 0),
      try1_call_reqs => try1_call_reqs(0 downto 0),
      try1_call_acks => try1_call_acks(0 downto 0),
      try1_call_tag => try1_call_tag(0 downto 0),
      try1_return_reqs => try1_return_reqs(0 downto 0),
      try1_return_acks => try1_return_acks(0 downto 0),
      try1_return_tag => try1_return_tag(0 downto 0),
      tag_in => try_tag_in,
      tag_out => try_tag_out-- 
    ); -- 
  -- module will be run forever 
  try_tag_in <= (others => '0');
  try_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => try_start_req, start_ack => try_start_ack,  fin_req => try_fin_req,  fin_ack => try_fin_ack);
  -- module try1
  -- call arbiter for module try1
  try1_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => try1_call_reqs,
      call_acks => try1_call_acks,
      return_reqs => try1_return_reqs,
      return_acks => try1_return_acks,
      call_tag  => try1_call_tag,
      return_tag  => try1_return_tag,
      call_mtag => try1_tag_in,
      return_mtag => try1_tag_out,
      call_mreq => try1_start_req,
      call_mack => try1_start_ack,
      return_mreq => try1_fin_req,
      return_mack => try1_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  try1_instance:try1-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => try1_start_req,
      start_ack => try1_start_ack,
      fin_req => try1_fin_req,
      fin_ack => try1_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(0 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(19 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(15 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(2 downto 0),
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(0 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(11 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(3 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(17 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(15 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(3 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(20 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(15 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(3 downto 0),
      memory_space_4_lr_req => memory_space_4_lr_req(0 downto 0),
      memory_space_4_lr_ack => memory_space_4_lr_ack(0 downto 0),
      memory_space_4_lr_addr => memory_space_4_lr_addr(3 downto 0),
      memory_space_4_lr_tag => memory_space_4_lr_tag(19 downto 0),
      memory_space_4_lc_req => memory_space_4_lc_req(0 downto 0),
      memory_space_4_lc_ack => memory_space_4_lc_ack(0 downto 0),
      memory_space_4_lc_data => memory_space_4_lc_data(15 downto 0),
      memory_space_4_lc_tag => memory_space_4_lc_tag(2 downto 0),
      memory_space_5_lr_req => memory_space_5_lr_req(0 downto 0),
      memory_space_5_lr_ack => memory_space_5_lr_ack(0 downto 0),
      memory_space_5_lr_addr => memory_space_5_lr_addr(10 downto 0),
      memory_space_5_lr_tag => memory_space_5_lr_tag(20 downto 0),
      memory_space_5_lc_req => memory_space_5_lc_req(0 downto 0),
      memory_space_5_lc_ack => memory_space_5_lc_ack(0 downto 0),
      memory_space_5_lc_data => memory_space_5_lc_data(15 downto 0),
      memory_space_5_lc_tag => memory_space_5_lc_tag(2 downto 0),
      memory_space_6_lr_req => memory_space_6_lr_req(0 downto 0),
      memory_space_6_lr_ack => memory_space_6_lr_ack(0 downto 0),
      memory_space_6_lr_addr => memory_space_6_lr_addr(0 downto 0),
      memory_space_6_lr_tag => memory_space_6_lr_tag(18 downto 0),
      memory_space_6_lc_req => memory_space_6_lc_req(0 downto 0),
      memory_space_6_lc_ack => memory_space_6_lc_ack(0 downto 0),
      memory_space_6_lc_data => memory_space_6_lc_data(0 downto 0),
      memory_space_6_lc_tag => memory_space_6_lc_tag(1 downto 0),
      memory_space_7_lr_req => memory_space_7_lr_req(0 downto 0),
      memory_space_7_lr_ack => memory_space_7_lr_ack(0 downto 0),
      memory_space_7_lr_addr => memory_space_7_lr_addr(0 downto 0),
      memory_space_7_lr_tag => memory_space_7_lr_tag(18 downto 0),
      memory_space_7_lc_req => memory_space_7_lc_req(0 downto 0),
      memory_space_7_lc_ack => memory_space_7_lc_ack(0 downto 0),
      memory_space_7_lc_data => memory_space_7_lc_data(15 downto 0),
      memory_space_7_lc_tag => memory_space_7_lc_tag(1 downto 0),
      memory_space_8_lr_req => memory_space_8_lr_req(0 downto 0),
      memory_space_8_lr_ack => memory_space_8_lr_ack(0 downto 0),
      memory_space_8_lr_addr => memory_space_8_lr_addr(0 downto 0),
      memory_space_8_lr_tag => memory_space_8_lr_tag(17 downto 0),
      memory_space_8_lc_req => memory_space_8_lc_req(0 downto 0),
      memory_space_8_lc_ack => memory_space_8_lc_ack(0 downto 0),
      memory_space_8_lc_data => memory_space_8_lc_data(3 downto 0),
      memory_space_8_lc_tag => memory_space_8_lc_tag(0 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(0 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(15 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(19 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(2 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(3 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(15 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(17 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(3 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(15 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(20 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(3 downto 0),
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(3 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(15 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(19 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(2 downto 0),
      memory_space_7_sr_req => memory_space_7_sr_req(0 downto 0),
      memory_space_7_sr_ack => memory_space_7_sr_ack(0 downto 0),
      memory_space_7_sr_addr => memory_space_7_sr_addr(0 downto 0),
      memory_space_7_sr_data => memory_space_7_sr_data(15 downto 0),
      memory_space_7_sr_tag => memory_space_7_sr_tag(18 downto 0),
      memory_space_7_sc_req => memory_space_7_sc_req(0 downto 0),
      memory_space_7_sc_ack => memory_space_7_sc_ack(0 downto 0),
      memory_space_7_sc_tag => memory_space_7_sc_tag(1 downto 0),
      acc_mem_pipe_write_req => acc_mem_pipe_write_req(0 downto 0),
      acc_mem_pipe_write_ack => acc_mem_pipe_write_ack(0 downto 0),
      acc_mem_pipe_write_data => acc_mem_pipe_write_data(15 downto 0),
      acc_mem_add_pipe_write_req => acc_mem_add_pipe_write_req(0 downto 0),
      acc_mem_add_pipe_write_ack => acc_mem_add_pipe_write_ack(0 downto 0),
      acc_mem_add_pipe_write_data => acc_mem_add_pipe_write_data(15 downto 0),
      accessMem_call_reqs => accessMem_call_reqs(2 downto 2),
      accessMem_call_acks => accessMem_call_acks(2 downto 2),
      accessMem_call_data => accessMem_call_data(86 downto 58),
      accessMem_call_tag => accessMem_call_tag(5 downto 4),
      accessMem_return_reqs => accessMem_return_reqs(2 downto 2),
      accessMem_return_acks => accessMem_return_acks(2 downto 2),
      accessMem_return_data => accessMem_return_data(191 downto 128),
      accessMem_return_tag => accessMem_return_tag(5 downto 4),
      accMemAccessDaemon_call_reqs => accMemAccessDaemon_call_reqs(0 downto 0),
      accMemAccessDaemon_call_acks => accMemAccessDaemon_call_acks(0 downto 0),
      accMemAccessDaemon_call_data => accMemAccessDaemon_call_data(31 downto 0),
      accMemAccessDaemon_call_tag => accMemAccessDaemon_call_tag(1 downto 0),
      accMemAccessDaemon_return_reqs => accMemAccessDaemon_return_reqs(0 downto 0),
      accMemAccessDaemon_return_acks => accMemAccessDaemon_return_acks(0 downto 0),
      accMemAccessDaemon_return_data => accMemAccessDaemon_return_data(63 downto 0),
      accMemAccessDaemon_return_tag => accMemAccessDaemon_return_tag(1 downto 0),
      accessMem_v_call_reqs => accessMem_v_call_reqs(0 downto 0),
      accessMem_v_call_acks => accessMem_v_call_acks(0 downto 0),
      accessMem_v_call_data => accessMem_v_call_data(28 downto 0),
      accessMem_v_call_tag => accessMem_v_call_tag(0 downto 0),
      accessMem_v_return_reqs => accessMem_v_return_reqs(0 downto 0),
      accessMem_v_return_acks => accessMem_v_return_acks(0 downto 0),
      accessMem_v_return_data => accessMem_v_return_data(63 downto 0),
      accessMem_v_return_tag => accessMem_v_return_tag(0 downto 0),
      tag_in => try1_tag_in,
      tag_out => try1_tag_out-- 
    ); -- 
  acc_mem_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe acc_mem",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => acc_mem_pipe_read_req,
      read_ack => acc_mem_pipe_read_ack,
      read_data => acc_mem_pipe_read_data,
      write_req => acc_mem_pipe_write_req,
      write_ack => acc_mem_pipe_write_ack,
      write_data => acc_mem_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  acc_mem_add_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe acc_mem_add",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => acc_mem_add_pipe_read_req,
      read_ack => acc_mem_add_pipe_read_ack,
      read_data => acc_mem_add_pipe_read_data,
      write_req => acc_mem_add_pipe_write_req,
      write_ack => acc_mem_add_pipe_write_ack,
      write_data => acc_mem_add_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => start_pipe_read_req,
      read_ack => start_pipe_read_ack,
      read_data => start_pipe_read_data,
      write_req => start_pipe_write_req,
      write_ack => start_pipe_write_ack,
      write_data => start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  status_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe status",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => status_pipe_read_req,
      read_ack => status_pipe_read_ack,
      read_data => status_pipe_read_data,
      write_req => status_pipe_write_req,
      write_ack => status_pipe_write_ack,
      write_data => status_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 2,
      num_stores => 1,
      addr_width => 1,
      data_width => 12,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 12
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 4,
      data_width => 16,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 4,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 1,
      num_stores => 1,
      addr_width => 4,
      data_width => 16,
      tag_width => 4,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 4,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_4: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_4",
      num_loads => 1,
      num_stores => 1,
      addr_width => 4,
      data_width => 16,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 4,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_4_lr_addr,
      lr_req_in => memory_space_4_lr_req,
      lr_ack_out => memory_space_4_lr_ack,
      lr_tag_in => memory_space_4_lr_tag,
      lc_req_in => memory_space_4_lc_req,
      lc_ack_out => memory_space_4_lc_ack,
      lc_data_out => memory_space_4_lc_data,
      lc_tag_out => memory_space_4_lc_tag,
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_5: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_5",
      num_loads => 3,
      num_stores => 2,
      addr_width => 11,
      data_width => 16,
      tag_width => 3,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 11,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_5_lr_addr,
      lr_req_in => memory_space_5_lr_req,
      lr_ack_out => memory_space_5_lr_ack,
      lr_tag_in => memory_space_5_lr_tag,
      lc_req_in => memory_space_5_lc_req,
      lc_ack_out => memory_space_5_lc_ack,
      lc_data_out => memory_space_5_lc_data,
      lc_tag_out => memory_space_5_lc_tag,
      sr_addr_in => memory_space_5_sr_addr,
      sr_data_in => memory_space_5_sr_data,
      sr_req_in => memory_space_5_sr_req,
      sr_ack_out => memory_space_5_sr_ack,
      sr_tag_in => memory_space_5_sr_tag,
      sc_req_in=> memory_space_5_sc_req,
      sc_ack_out => memory_space_5_sc_ack,
      sc_tag_out => memory_space_5_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_6: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_6",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 1,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 1
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_6_lr_addr,
      lr_req_in => memory_space_6_lr_req,
      lr_ack_out => memory_space_6_lr_ack,
      lr_tag_in => memory_space_6_lr_tag,
      lc_req_in => memory_space_6_lc_req,
      lc_ack_out => memory_space_6_lc_ack,
      lc_data_out => memory_space_6_lc_data,
      lc_tag_out => memory_space_6_lc_tag,
      sr_addr_in => memory_space_6_sr_addr,
      sr_data_in => memory_space_6_sr_data,
      sr_req_in => memory_space_6_sr_req,
      sr_ack_out => memory_space_6_sr_ack,
      sr_tag_in => memory_space_6_sr_tag,
      sc_req_in=> memory_space_6_sc_req,
      sc_ack_out => memory_space_6_sc_ack,
      sc_tag_out => memory_space_6_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_7: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_7",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_7_lr_addr,
      lr_req_in => memory_space_7_lr_req,
      lr_ack_out => memory_space_7_lr_ack,
      lr_tag_in => memory_space_7_lr_tag,
      lc_req_in => memory_space_7_lc_req,
      lc_ack_out => memory_space_7_lc_ack,
      lc_data_out => memory_space_7_lc_data,
      lc_tag_out => memory_space_7_lc_tag,
      sr_addr_in => memory_space_7_sr_addr,
      sr_data_in => memory_space_7_sr_data,
      sr_req_in => memory_space_7_sr_req,
      sr_ack_out => memory_space_7_sr_ack,
      sr_tag_in => memory_space_7_sr_tag,
      sc_req_in=> memory_space_7_sc_req,
      sc_ack_out => memory_space_7_sc_ack,
      sc_tag_out => memory_space_7_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_8: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_8",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 4,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 4
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_8_lr_addr,
      lr_req_in => memory_space_8_lr_req,
      lr_ack_out => memory_space_8_lr_ack,
      lr_tag_in => memory_space_8_lr_tag,
      lc_req_in => memory_space_8_lc_req,
      lc_ack_out => memory_space_8_lc_ack,
      lc_data_out => memory_space_8_lc_data,
      lc_tag_out => memory_space_8_lc_tag,
      sr_addr_in => memory_space_8_sr_addr,
      sr_data_in => memory_space_8_sr_data,
      sr_req_in => memory_space_8_sr_req,
      sr_ack_out => memory_space_8_sr_ack,
      sr_tag_in => memory_space_8_sr_tag,
      sc_req_in=> memory_space_8_sc_req,
      sc_ack_out => memory_space_8_sc_ack,
      sc_tag_out => memory_space_8_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
