-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity accessMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    read_write_bar : in  std_logic_vector(0 downto 0);
    addr : in  std_logic_vector(7 downto 0);
    write_data : in  std_logic_vector(31 downto 0);
    read_data : out  std_logic_vector(31 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(7 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(7 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessMem;
architecture accessMem_arch of accessMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 41)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal read_write_bar_buffer :  std_logic_vector(0 downto 0);
  signal read_write_bar_update_enable: Boolean;
  signal addr_buffer :  std_logic_vector(7 downto 0);
  signal addr_update_enable: Boolean;
  signal write_data_buffer :  std_logic_vector(31 downto 0);
  signal write_data_update_enable: Boolean;
  -- output port buffer signals
  signal read_data_buffer :  std_logic_vector(31 downto 0);
  signal read_data_update_enable: Boolean;
  signal accessMem_CP_0_start: Boolean;
  signal accessMem_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_19_store_0_req_1 : boolean;
  signal array_obj_ref_19_store_0_ack_1 : boolean;
  signal array_obj_ref_19_store_0_req_0 : boolean;
  signal array_obj_ref_19_store_0_ack_0 : boolean;
  signal array_obj_ref_25_load_0_req_0 : boolean;
  signal array_obj_ref_25_load_0_ack_0 : boolean;
  signal array_obj_ref_25_load_0_req_1 : boolean;
  signal array_obj_ref_25_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessMem_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 41) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= read_write_bar;
  read_write_bar_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(8 downto 1) <= addr;
  addr_buffer <= in_buffer_data_out(8 downto 1);
  in_buffer_data_in(40 downto 9) <= write_data;
  write_data_buffer <= in_buffer_data_out(40 downto 9);
  in_buffer_data_in(tag_length + 40 downto 41) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 40 downto 41);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 7,2 => 7,3 => 1,4 => 7);
    constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 7);
    constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 5); -- 
  begin -- 
    preds <= read_write_bar_update_enable & addr_update_enable & write_data_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessMem_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= read_data_buffer;
  read_data <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMem_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  read_data_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 28) := "read_data_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_read_data_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => read_data_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 7,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessMem_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMem_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessMem_CP_0: Block -- control-path 
    signal accessMem_CP_0_elements: BooleanArray(21 downto 0);
    -- 
  begin -- 
    accessMem_CP_0_elements(0) <= accessMem_CP_0_start;
    accessMem_CP_0_symbol <= accessMem_CP_0_elements(21);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	10 
    -- CP-element group 1: 	6 
    -- CP-element group 1:  members (53) 
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/$entry
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_index_computed_0
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_index_resize_0/$entry
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_index_resize_0/$exit
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_index_resize_0/index_resize_req
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_index_resize_0/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_index_scale_0/$entry
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_index_scale_0/$exit
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_index_scale_0/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_index_scale_0/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_final_index_sum_regn/$entry
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_final_index_sum_regn/$exit
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_word_address_calculated
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_root_address_calculated
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_offset_calculated
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_index_resized_0
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_index_scaled_0
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_final_index_sum_regn/req
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_final_index_sum_regn/ack
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_base_plus_offset/$entry
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_base_plus_offset/$exit
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_base_plus_offset/sum_rename_req
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_base_plus_offset/sum_rename_ack
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_word_addrgen/$entry
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_word_addrgen/$exit
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_word_addrgen/root_register_req
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_word_addrgen/root_register_ack
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_word_address_calculated
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_root_address_calculated
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_offset_calculated
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_index_resized_0
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_index_scaled_0
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_index_computed_0
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_index_resize_0/$entry
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_index_resize_0/$exit
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_index_resize_0/index_resize_req
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_index_resize_0/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_index_scale_0/$entry
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_index_scale_0/$exit
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_index_scale_0/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_index_scale_0/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_final_index_sum_regn/$entry
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_final_index_sum_regn/$exit
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_final_index_sum_regn/req
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_final_index_sum_regn/ack
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_base_plus_offset/$entry
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_base_plus_offset/$exit
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_base_plus_offset/sum_rename_req
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_base_plus_offset/sum_rename_ack
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_word_addrgen/$entry
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_word_addrgen/$exit
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_word_addrgen/root_register_req
      -- CP-element group 1: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_word_addrgen/root_register_ack
      -- 
    accessMem_CP_0_elements(1) <= accessMem_CP_0_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	12 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	17 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_21_to_assign_stmt_26/read_write_bar_update_enable
      -- CP-element group 2: 	 assign_stmt_21_to_assign_stmt_26/read_write_bar_update_enable_out
      -- 
    accessMem_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "accessMem_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(8) & accessMem_CP_0_elements(12);
      gj_accessMem_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	8 
    -- CP-element group 3: 	12 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	18 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_21_to_assign_stmt_26/addr_update_enable
      -- CP-element group 3: 	 assign_stmt_21_to_assign_stmt_26/addr_update_enable_out
      -- 
    accessMem_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "accessMem_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(8) & accessMem_CP_0_elements(12);
      gj_accessMem_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	8 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	19 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_21_to_assign_stmt_26/write_data_update_enable_out
      -- CP-element group 4: 	 assign_stmt_21_to_assign_stmt_26/write_data_update_enable
      -- 
    accessMem_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "accessMem_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMem_CP_0_elements(8);
      gj_accessMem_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	20 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	11 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_21_to_assign_stmt_26/read_data_update_enable
      -- CP-element group 5: 	 assign_stmt_21_to_assign_stmt_26/read_data_update_enable_in
      -- 
    accessMem_CP_0_elements(5) <= accessMem_CP_0_elements(20);
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	1 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	8 
    -- CP-element group 6: 	15 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_sample_start_
      -- CP-element group 6: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_Sample/$entry
      -- CP-element group 6: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_Sample/array_obj_ref_19_Split/$entry
      -- CP-element group 6: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_Sample/array_obj_ref_19_Split/$exit
      -- CP-element group 6: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_Sample/array_obj_ref_19_Split/split_req
      -- CP-element group 6: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_Sample/array_obj_ref_19_Split/split_ack
      -- CP-element group 6: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_Sample/word_access_start/$entry
      -- CP-element group 6: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_Sample/word_access_start/word_0/$entry
      -- CP-element group 6: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_Sample/word_access_start/word_0/rr
      -- 
    rr_63_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_63_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(6), ack => array_obj_ref_19_store_0_req_0); -- 
    accessMem_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 28) := "accessMem_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(8) & accessMem_CP_0_elements(15);
      gj_accessMem_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: marked-predecessors 
    -- CP-element group 7: 	9 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	9 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_Update/word_access_complete/word_0/$entry
      -- CP-element group 7: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_Update/word_access_complete/word_0/cr
      -- CP-element group 7: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_update_start_
      -- CP-element group 7: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_Update/$entry
      -- CP-element group 7: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_Update/word_access_complete/$entry
      -- 
    cr_74_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_74_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(7), ack => array_obj_ref_19_store_0_req_1); -- 
    accessMem_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "accessMem_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMem_CP_0_elements(9);
      gj_accessMem_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	14 
    -- CP-element group 8: 	15 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	3 
    -- CP-element group 8: 	4 
    -- CP-element group 8: 	2 
    -- CP-element group 8: 	6 
    -- CP-element group 8:  members (5) 
      -- CP-element group 8: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_sample_completed_
      -- CP-element group 8: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_Sample/$exit
      -- CP-element group 8: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_Sample/word_access_start/$exit
      -- CP-element group 8: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_Sample/word_access_start/word_0/$exit
      -- CP-element group 8: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_Sample/word_access_start/word_0/ra
      -- 
    ra_64_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_19_store_0_ack_0, ack => accessMem_CP_0_elements(8)); -- 
    -- CP-element group 9:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	7 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	16 
    -- CP-element group 9: marked-successors 
    -- CP-element group 9: 	7 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_Update/word_access_complete/word_0/$exit
      -- CP-element group 9: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_Update/word_access_complete/word_0/ca
      -- CP-element group 9: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_update_completed_
      -- CP-element group 9: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_Update/$exit
      -- CP-element group 9: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_Update/word_access_complete/$exit
      -- 
    ca_75_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_19_store_0_ack_1, ack => accessMem_CP_0_elements(9)); -- 
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	1 
    -- CP-element group 10: 	14 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (5) 
      -- CP-element group 10: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_sample_start_
      -- CP-element group 10: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_Sample/word_access_start/$entry
      -- CP-element group 10: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_Sample/word_access_start/word_0/$entry
      -- CP-element group 10: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_Sample/word_access_start/word_0/rr
      -- 
    rr_121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(10), ack => array_obj_ref_25_load_0_req_0); -- 
    accessMem_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(14) & accessMem_CP_0_elements(12);
      gj_accessMem_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	5 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	13 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_update_start_
      -- CP-element group 11: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_Update/$entry
      -- CP-element group 11: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_Update/word_access_complete/$entry
      -- CP-element group 11: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_Update/word_access_complete/word_0/$entry
      -- CP-element group 11: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_Update/word_access_complete/word_0/cr
      -- 
    cr_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(11), ack => array_obj_ref_25_load_0_req_1); -- 
    accessMem_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(5) & accessMem_CP_0_elements(13);
      gj_accessMem_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: 	3 
    -- CP-element group 12: 	2 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_sample_completed_
      -- CP-element group 12: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_Sample/$exit
      -- CP-element group 12: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_Sample/word_access_start/$exit
      -- CP-element group 12: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_Sample/word_access_start/word_0/$exit
      -- CP-element group 12: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_Sample/word_access_start/word_0/ra
      -- 
    ra_122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_25_load_0_ack_0, ack => accessMem_CP_0_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	11 
    -- CP-element group 13:  members (9) 
      -- CP-element group 13: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_update_completed_
      -- CP-element group 13: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_Update/$exit
      -- CP-element group 13: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_Update/word_access_complete/$exit
      -- CP-element group 13: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_Update/word_access_complete/word_0/$exit
      -- CP-element group 13: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_Update/word_access_complete/word_0/ca
      -- CP-element group 13: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_Update/array_obj_ref_25_Merge/$entry
      -- CP-element group 13: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_Update/array_obj_ref_25_Merge/$exit
      -- CP-element group 13: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_Update/array_obj_ref_25_Merge/merge_req
      -- CP-element group 13: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_25_Update/array_obj_ref_25_Merge/merge_ack
      -- 
    ca_133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_25_load_0_ack_1, ack => accessMem_CP_0_elements(13)); -- 
    -- CP-element group 14:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	8 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 assign_stmt_21_to_assign_stmt_26/array_obj_ref_19_array_obj_ref_25_delay
      -- 
    -- Element group accessMem_CP_0_elements(14) is a control-delay.
    cp_element_14_delay: control_delay_element  generic map(name => " 14_delay", delay_value => 1)  port map(req => accessMem_CP_0_elements(8), ack => accessMem_CP_0_elements(14), clk => clk, reset =>reset);
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	8 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	6 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 assign_stmt_21_to_assign_stmt_26/ring_reenable_memory_space_0
      -- 
    accessMem_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(8) & accessMem_CP_0_elements(12);
      gj_accessMem_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: 	9 
    -- CP-element group 16: 	13 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	21 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 assign_stmt_21_to_assign_stmt_26/$exit
      -- 
    accessMem_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(15) & accessMem_CP_0_elements(9) & accessMem_CP_0_elements(13);
      gj_accessMem_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 read_write_bar_update_enable
      -- 
    accessMem_CP_0_elements(17) <= accessMem_CP_0_elements(2);
    -- CP-element group 18:  place  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	3 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 addr_update_enable
      -- 
    accessMem_CP_0_elements(18) <= accessMem_CP_0_elements(3);
    -- CP-element group 19:  place  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	4 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 write_data_update_enable
      -- 
    accessMem_CP_0_elements(19) <= accessMem_CP_0_elements(4);
    -- CP-element group 20:  place  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	5 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 read_data_update_enable
      -- 
    -- CP-element group 21:  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	16 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 $exit
      -- 
    accessMem_CP_0_elements(21) <= accessMem_CP_0_elements(16);
    --  hookup: inputs to control-path 
    accessMem_CP_0_elements(20) <= read_data_update_enable;
    -- hookup: output from control-path 
    read_write_bar_update_enable <= accessMem_CP_0_elements(17);
    addr_update_enable <= accessMem_CP_0_elements(18);
    write_data_update_enable <= accessMem_CP_0_elements(19);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_addr_18_resized : std_logic_vector(7 downto 0);
    signal R_addr_18_scaled : std_logic_vector(7 downto 0);
    signal R_addr_24_resized : std_logic_vector(7 downto 0);
    signal R_addr_24_scaled : std_logic_vector(7 downto 0);
    signal array_obj_ref_19_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_19_final_offset : std_logic_vector(7 downto 0);
    signal array_obj_ref_19_offset_scale_factor_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_19_resized_base_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_19_root_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_19_word_address_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_19_word_offset_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_25_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_25_final_offset : std_logic_vector(7 downto 0);
    signal array_obj_ref_25_offset_scale_factor_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_25_resized_base_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_25_root_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_25_word_address_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_25_word_offset_0 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_19_offset_scale_factor_0 <= "00000001";
    array_obj_ref_19_resized_base_address <= "00000000";
    array_obj_ref_19_word_offset_0 <= "00000000";
    array_obj_ref_25_offset_scale_factor_0 <= "00000001";
    array_obj_ref_25_resized_base_address <= "00000000";
    array_obj_ref_25_word_offset_0 <= "00000000";
    -- equivalence array_obj_ref_19_addr_0
    process(array_obj_ref_19_root_address) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_19_root_address;
      ov(7 downto 0) := iv;
      array_obj_ref_19_word_address_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_19_gather_scatter
    process(write_data_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := write_data_buffer;
      ov(31 downto 0) := iv;
      array_obj_ref_19_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_19_index_0_rename
    process(R_addr_18_resized) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_18_resized;
      ov(7 downto 0) := iv;
      R_addr_18_scaled <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_19_index_0_resize
    process(addr_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_buffer;
      ov(7 downto 0) := iv;
      R_addr_18_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_19_index_offset
    process(R_addr_18_scaled) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_18_scaled;
      ov(7 downto 0) := iv;
      array_obj_ref_19_final_offset <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_19_root_address_inst
    process(array_obj_ref_19_final_offset) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_19_final_offset;
      ov(7 downto 0) := iv;
      array_obj_ref_19_root_address <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_25_addr_0
    process(array_obj_ref_25_root_address) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_25_root_address;
      ov(7 downto 0) := iv;
      array_obj_ref_25_word_address_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_25_gather_scatter
    process(array_obj_ref_25_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_25_data_0;
      ov(31 downto 0) := iv;
      read_data_buffer <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_25_index_0_rename
    process(R_addr_24_resized) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_24_resized;
      ov(7 downto 0) := iv;
      R_addr_24_scaled <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_25_index_0_resize
    process(addr_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_buffer;
      ov(7 downto 0) := iv;
      R_addr_24_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_25_index_offset
    process(R_addr_24_scaled) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_24_scaled;
      ov(7 downto 0) := iv;
      array_obj_ref_25_final_offset <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_25_root_address_inst
    process(array_obj_ref_25_final_offset) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_25_final_offset;
      ov(7 downto 0) := iv;
      array_obj_ref_25_root_address <= ov(7 downto 0);
      --
    end process;
    -- shared load operator group (0) : array_obj_ref_25_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_25_load_0_req_0;
      array_obj_ref_25_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_25_load_0_req_1;
      array_obj_ref_25_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_write_bar_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_25_word_address_0;
      array_obj_ref_25_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 8,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(7 downto 0),
          mtag => memory_space_0_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : array_obj_ref_19_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(7 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 7);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_19_store_0_req_0;
      array_obj_ref_19_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_19_store_0_req_1;
      array_obj_ref_19_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_write_bar_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_19_word_address_0;
      data_in <= array_obj_ref_19_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 8,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(7 downto 0),
          mdata => memory_space_0_sr_data(31 downto 0),
          mtag => memory_space_0_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end accessMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity accessreg is -- 
  generic (tag_length : integer); 
  port ( -- 
    read_write_bar : in  std_logic_vector(0 downto 0);
    addr : in  std_logic_vector(7 downto 0);
    write_data : in  std_logic_vector(31 downto 0);
    read_data : out  std_logic_vector(31 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(7 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(7 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessreg;
architecture accessreg_arch of accessreg is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 41)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal read_write_bar_buffer :  std_logic_vector(0 downto 0);
  signal read_write_bar_update_enable: Boolean;
  signal addr_buffer :  std_logic_vector(7 downto 0);
  signal addr_update_enable: Boolean;
  signal write_data_buffer :  std_logic_vector(31 downto 0);
  signal write_data_update_enable: Boolean;
  -- output port buffer signals
  signal read_data_buffer :  std_logic_vector(31 downto 0);
  signal read_data_update_enable: Boolean;
  signal accessreg_CP_145_start: Boolean;
  signal accessreg_CP_145_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_35_store_0_ack_1 : boolean;
  signal array_obj_ref_35_store_0_req_0 : boolean;
  signal array_obj_ref_35_store_0_ack_0 : boolean;
  signal array_obj_ref_35_store_0_req_1 : boolean;
  signal array_obj_ref_41_load_0_req_0 : boolean;
  signal array_obj_ref_41_load_0_ack_0 : boolean;
  signal array_obj_ref_41_load_0_req_1 : boolean;
  signal array_obj_ref_41_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessreg_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 41) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= read_write_bar;
  read_write_bar_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(8 downto 1) <= addr;
  addr_buffer <= in_buffer_data_out(8 downto 1);
  in_buffer_data_in(40 downto 9) <= write_data;
  write_data_buffer <= in_buffer_data_out(40 downto 9);
  in_buffer_data_in(tag_length + 40 downto 41) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 40 downto 41);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 7,2 => 7,3 => 1,4 => 7);
    constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 7);
    constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 5); -- 
  begin -- 
    preds <= read_write_bar_update_enable & addr_update_enable & write_data_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessreg_CP_145_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessreg_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= read_data_buffer;
  read_data <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessreg_CP_145_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  read_data_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 28) := "read_data_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_read_data_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => read_data_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 7,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessreg_CP_145_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessreg_CP_145_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessreg_CP_145: Block -- control-path 
    signal accessreg_CP_145_elements: BooleanArray(21 downto 0);
    -- 
  begin -- 
    accessreg_CP_145_elements(0) <= accessreg_CP_145_start;
    accessreg_CP_145_symbol <= accessreg_CP_145_elements(21);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	10 
    -- CP-element group 1: 	6 
    -- CP-element group 1:  members (53) 
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/$entry
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_word_address_calculated
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_root_address_calculated
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_offset_calculated
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_index_resized_0
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_index_scaled_0
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_index_computed_0
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_index_resize_0/$entry
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_index_resize_0/$exit
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_index_resize_0/index_resize_req
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_index_resize_0/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_index_scale_0/$entry
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_index_scale_0/$exit
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_index_scale_0/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_index_scale_0/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_final_index_sum_regn/$entry
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_final_index_sum_regn/$exit
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_final_index_sum_regn/req
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_final_index_sum_regn/ack
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_base_plus_offset/$entry
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_base_plus_offset/$exit
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_base_plus_offset/sum_rename_req
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_base_plus_offset/sum_rename_ack
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_word_addrgen/$entry
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_word_addrgen/$exit
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_word_addrgen/root_register_req
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_word_addrgen/root_register_ack
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_word_address_calculated
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_root_address_calculated
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_offset_calculated
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_index_resized_0
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_index_scaled_0
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_index_computed_0
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_index_resize_0/$entry
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_index_resize_0/$exit
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_index_resize_0/index_resize_req
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_index_resize_0/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_index_scale_0/$entry
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_index_scale_0/$exit
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_index_scale_0/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_index_scale_0/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_final_index_sum_regn/$entry
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_final_index_sum_regn/$exit
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_final_index_sum_regn/req
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_final_index_sum_regn/ack
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_base_plus_offset/$entry
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_base_plus_offset/$exit
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_base_plus_offset/sum_rename_req
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_base_plus_offset/sum_rename_ack
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_word_addrgen/$entry
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_word_addrgen/$exit
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_word_addrgen/root_register_req
      -- CP-element group 1: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_word_addrgen/root_register_ack
      -- 
    accessreg_CP_145_elements(1) <= accessreg_CP_145_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	8 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	17 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_37_to_assign_stmt_42/read_write_bar_update_enable
      -- CP-element group 2: 	 assign_stmt_37_to_assign_stmt_42/read_write_bar_update_enable_out
      -- 
    accessreg_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "accessreg_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessreg_CP_145_elements(12) & accessreg_CP_145_elements(8);
      gj_accessreg_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessreg_CP_145_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	12 
    -- CP-element group 3: 	8 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	18 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_37_to_assign_stmt_42/addr_update_enable
      -- CP-element group 3: 	 assign_stmt_37_to_assign_stmt_42/addr_update_enable_out
      -- 
    accessreg_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "accessreg_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessreg_CP_145_elements(12) & accessreg_CP_145_elements(8);
      gj_accessreg_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessreg_CP_145_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	8 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	19 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_37_to_assign_stmt_42/write_data_update_enable
      -- CP-element group 4: 	 assign_stmt_37_to_assign_stmt_42/write_data_update_enable_out
      -- 
    accessreg_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "accessreg_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessreg_CP_145_elements(8);
      gj_accessreg_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessreg_CP_145_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	20 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	11 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_37_to_assign_stmt_42/read_data_update_enable
      -- CP-element group 5: 	 assign_stmt_37_to_assign_stmt_42/read_data_update_enable_in
      -- 
    accessreg_CP_145_elements(5) <= accessreg_CP_145_elements(20);
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	1 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	15 
    -- CP-element group 6: 	8 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_sample_start_
      -- CP-element group 6: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_Sample/$entry
      -- CP-element group 6: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_Sample/array_obj_ref_35_Split/$entry
      -- CP-element group 6: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_Sample/array_obj_ref_35_Split/$exit
      -- CP-element group 6: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_Sample/array_obj_ref_35_Split/split_req
      -- CP-element group 6: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_Sample/array_obj_ref_35_Split/split_ack
      -- CP-element group 6: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_Sample/word_access_start/$entry
      -- CP-element group 6: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_Sample/word_access_start/word_0/$entry
      -- CP-element group 6: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_Sample/word_access_start/word_0/rr
      -- 
    rr_208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessreg_CP_145_elements(6), ack => array_obj_ref_35_store_0_req_0); -- 
    accessreg_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 28) := "accessreg_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessreg_CP_145_elements(1) & accessreg_CP_145_elements(15) & accessreg_CP_145_elements(8);
      gj_accessreg_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessreg_CP_145_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: marked-predecessors 
    -- CP-element group 7: 	9 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	9 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_update_start_
      -- CP-element group 7: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_Update/$entry
      -- CP-element group 7: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_Update/word_access_complete/$entry
      -- CP-element group 7: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_Update/word_access_complete/word_0/$entry
      -- CP-element group 7: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_Update/word_access_complete/word_0/cr
      -- 
    cr_219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessreg_CP_145_elements(7), ack => array_obj_ref_35_store_0_req_1); -- 
    accessreg_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "accessreg_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessreg_CP_145_elements(9);
      gj_accessreg_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessreg_CP_145_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	14 
    -- CP-element group 8: 	15 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	4 
    -- CP-element group 8: 	2 
    -- CP-element group 8: 	3 
    -- CP-element group 8: 	6 
    -- CP-element group 8:  members (5) 
      -- CP-element group 8: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_sample_completed_
      -- CP-element group 8: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_Sample/$exit
      -- CP-element group 8: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_Sample/word_access_start/$exit
      -- CP-element group 8: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_Sample/word_access_start/word_0/$exit
      -- CP-element group 8: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_Sample/word_access_start/word_0/ra
      -- 
    ra_209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_35_store_0_ack_0, ack => accessreg_CP_145_elements(8)); -- 
    -- CP-element group 9:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	7 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	16 
    -- CP-element group 9: marked-successors 
    -- CP-element group 9: 	7 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_Update/word_access_complete/word_0/ca
      -- CP-element group 9: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_update_completed_
      -- CP-element group 9: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_Update/$exit
      -- CP-element group 9: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_Update/word_access_complete/$exit
      -- CP-element group 9: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_Update/word_access_complete/word_0/$exit
      -- 
    ca_220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_35_store_0_ack_1, ack => accessreg_CP_145_elements(9)); -- 
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	1 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (5) 
      -- CP-element group 10: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_sample_start_
      -- CP-element group 10: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_Sample/word_access_start/$entry
      -- CP-element group 10: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_Sample/word_access_start/word_0/$entry
      -- CP-element group 10: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_Sample/word_access_start/word_0/rr
      -- 
    rr_266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessreg_CP_145_elements(10), ack => array_obj_ref_41_load_0_req_0); -- 
    accessreg_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "accessreg_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessreg_CP_145_elements(14) & accessreg_CP_145_elements(1) & accessreg_CP_145_elements(12);
      gj_accessreg_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessreg_CP_145_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	5 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	13 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_update_start_
      -- CP-element group 11: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_Update/$entry
      -- CP-element group 11: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_Update/word_access_complete/$entry
      -- CP-element group 11: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_Update/word_access_complete/word_0/$entry
      -- CP-element group 11: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_Update/word_access_complete/word_0/cr
      -- 
    cr_277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessreg_CP_145_elements(11), ack => array_obj_ref_41_load_0_req_1); -- 
    accessreg_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessreg_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessreg_CP_145_elements(5) & accessreg_CP_145_elements(13);
      gj_accessreg_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessreg_CP_145_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: 	2 
    -- CP-element group 12: 	3 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_sample_completed_
      -- CP-element group 12: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_Sample/$exit
      -- CP-element group 12: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_Sample/word_access_start/$exit
      -- CP-element group 12: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_Sample/word_access_start/word_0/$exit
      -- CP-element group 12: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_Sample/word_access_start/word_0/ra
      -- 
    ra_267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_41_load_0_ack_0, ack => accessreg_CP_145_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	11 
    -- CP-element group 13:  members (9) 
      -- CP-element group 13: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_update_completed_
      -- CP-element group 13: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_Update/$exit
      -- CP-element group 13: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_Update/word_access_complete/$exit
      -- CP-element group 13: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_Update/word_access_complete/word_0/$exit
      -- CP-element group 13: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_Update/word_access_complete/word_0/ca
      -- CP-element group 13: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_Update/array_obj_ref_41_Merge/$entry
      -- CP-element group 13: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_Update/array_obj_ref_41_Merge/$exit
      -- CP-element group 13: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_Update/array_obj_ref_41_Merge/merge_req
      -- CP-element group 13: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_41_Update/array_obj_ref_41_Merge/merge_ack
      -- 
    ca_278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_41_load_0_ack_1, ack => accessreg_CP_145_elements(13)); -- 
    -- CP-element group 14:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	8 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 assign_stmt_37_to_assign_stmt_42/array_obj_ref_35_array_obj_ref_41_delay
      -- 
    -- Element group accessreg_CP_145_elements(14) is a control-delay.
    cp_element_14_delay: control_delay_element  generic map(name => " 14_delay", delay_value => 1)  port map(req => accessreg_CP_145_elements(8), ack => accessreg_CP_145_elements(14), clk => clk, reset =>reset);
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: 	8 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	6 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 assign_stmt_37_to_assign_stmt_42/ring_reenable_memory_space_2
      -- 
    accessreg_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessreg_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessreg_CP_145_elements(12) & accessreg_CP_145_elements(8);
      gj_accessreg_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessreg_CP_145_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: 	13 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	21 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 assign_stmt_37_to_assign_stmt_42/$exit
      -- 
    accessreg_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "accessreg_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessreg_CP_145_elements(9) & accessreg_CP_145_elements(13) & accessreg_CP_145_elements(15);
      gj_accessreg_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessreg_CP_145_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 read_write_bar_update_enable
      -- 
    accessreg_CP_145_elements(17) <= accessreg_CP_145_elements(2);
    -- CP-element group 18:  place  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	3 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 addr_update_enable
      -- 
    accessreg_CP_145_elements(18) <= accessreg_CP_145_elements(3);
    -- CP-element group 19:  place  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	4 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 write_data_update_enable
      -- 
    accessreg_CP_145_elements(19) <= accessreg_CP_145_elements(4);
    -- CP-element group 20:  place  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	5 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 read_data_update_enable
      -- 
    -- CP-element group 21:  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	16 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 $exit
      -- 
    accessreg_CP_145_elements(21) <= accessreg_CP_145_elements(16);
    --  hookup: inputs to control-path 
    accessreg_CP_145_elements(20) <= read_data_update_enable;
    -- hookup: output from control-path 
    read_write_bar_update_enable <= accessreg_CP_145_elements(17);
    addr_update_enable <= accessreg_CP_145_elements(18);
    write_data_update_enable <= accessreg_CP_145_elements(19);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_addr_34_resized : std_logic_vector(7 downto 0);
    signal R_addr_34_scaled : std_logic_vector(7 downto 0);
    signal R_addr_40_resized : std_logic_vector(7 downto 0);
    signal R_addr_40_scaled : std_logic_vector(7 downto 0);
    signal array_obj_ref_35_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_35_final_offset : std_logic_vector(7 downto 0);
    signal array_obj_ref_35_offset_scale_factor_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_35_resized_base_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_35_root_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_35_word_address_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_35_word_offset_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_41_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_41_final_offset : std_logic_vector(7 downto 0);
    signal array_obj_ref_41_offset_scale_factor_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_41_resized_base_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_41_root_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_41_word_address_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_41_word_offset_0 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_35_offset_scale_factor_0 <= "00000001";
    array_obj_ref_35_resized_base_address <= "00000000";
    array_obj_ref_35_word_offset_0 <= "00000000";
    array_obj_ref_41_offset_scale_factor_0 <= "00000001";
    array_obj_ref_41_resized_base_address <= "00000000";
    array_obj_ref_41_word_offset_0 <= "00000000";
    -- equivalence array_obj_ref_35_addr_0
    process(array_obj_ref_35_root_address) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_35_root_address;
      ov(7 downto 0) := iv;
      array_obj_ref_35_word_address_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_35_gather_scatter
    process(write_data_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := write_data_buffer;
      ov(31 downto 0) := iv;
      array_obj_ref_35_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_35_index_0_rename
    process(R_addr_34_resized) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_34_resized;
      ov(7 downto 0) := iv;
      R_addr_34_scaled <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_35_index_0_resize
    process(addr_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_buffer;
      ov(7 downto 0) := iv;
      R_addr_34_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_35_index_offset
    process(R_addr_34_scaled) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_34_scaled;
      ov(7 downto 0) := iv;
      array_obj_ref_35_final_offset <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_35_root_address_inst
    process(array_obj_ref_35_final_offset) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_35_final_offset;
      ov(7 downto 0) := iv;
      array_obj_ref_35_root_address <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_41_addr_0
    process(array_obj_ref_41_root_address) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_41_root_address;
      ov(7 downto 0) := iv;
      array_obj_ref_41_word_address_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_41_gather_scatter
    process(array_obj_ref_41_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_41_data_0;
      ov(31 downto 0) := iv;
      read_data_buffer <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_41_index_0_rename
    process(R_addr_40_resized) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_40_resized;
      ov(7 downto 0) := iv;
      R_addr_40_scaled <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_41_index_0_resize
    process(addr_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_buffer;
      ov(7 downto 0) := iv;
      R_addr_40_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_41_index_offset
    process(R_addr_40_scaled) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_40_scaled;
      ov(7 downto 0) := iv;
      array_obj_ref_41_final_offset <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_41_root_address_inst
    process(array_obj_ref_41_final_offset) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_41_final_offset;
      ov(7 downto 0) := iv;
      array_obj_ref_41_root_address <= ov(7 downto 0);
      --
    end process;
    -- shared load operator group (0) : array_obj_ref_41_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_41_load_0_req_0;
      array_obj_ref_41_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_41_load_0_req_1;
      array_obj_ref_41_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_write_bar_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_41_word_address_0;
      array_obj_ref_41_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 8,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(7 downto 0),
          mtag => memory_space_2_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : array_obj_ref_35_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(7 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 7);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_35_store_0_req_0;
      array_obj_ref_35_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_35_store_0_req_1;
      array_obj_ref_35_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_write_bar_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_35_word_address_0;
      data_in <= array_obj_ref_35_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 8,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(7 downto 0),
          mdata => memory_space_2_sr_data(31 downto 0),
          mtag => memory_space_2_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end accessreg_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity add is -- 
  generic (tag_length : integer); 
  port ( -- 
    rs1_data : in  std_logic_vector(31 downto 0);
    rs2_data : in  std_logic_vector(31 downto 0);
    rd : in  std_logic_vector(7 downto 0);
    pc : in  std_logic_vector(7 downto 0);
    next_pc : out  std_logic_vector(7 downto 0);
    accessreg_call_reqs : out  std_logic_vector(0 downto 0);
    accessreg_call_acks : in   std_logic_vector(0 downto 0);
    accessreg_call_data : out  std_logic_vector(40 downto 0);
    accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
    accessreg_return_reqs : out  std_logic_vector(0 downto 0);
    accessreg_return_acks : in   std_logic_vector(0 downto 0);
    accessreg_return_data : in   std_logic_vector(31 downto 0);
    accessreg_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity add;
architecture add_arch of add is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 80)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rs1_data_buffer :  std_logic_vector(31 downto 0);
  signal rs1_data_update_enable: Boolean;
  signal rs2_data_buffer :  std_logic_vector(31 downto 0);
  signal rs2_data_update_enable: Boolean;
  signal rd_buffer :  std_logic_vector(7 downto 0);
  signal rd_update_enable: Boolean;
  signal pc_buffer :  std_logic_vector(7 downto 0);
  signal pc_update_enable: Boolean;
  -- output port buffer signals
  signal next_pc_buffer :  std_logic_vector(7 downto 0);
  signal next_pc_update_enable: Boolean;
  signal add_CP_290_start: Boolean;
  signal add_CP_290_symbol: Boolean;
  -- volatile/operator module components. 
  component accessreg is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(7 downto 0);
      write_data : in  std_logic_vector(31 downto 0);
      read_data : out  std_logic_vector(31 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal ADD_u32_u32_53_inst_req_0 : boolean;
  signal ADD_u32_u32_53_inst_ack_0 : boolean;
  signal ADD_u32_u32_53_inst_req_1 : boolean;
  signal ADD_u32_u32_53_inst_ack_1 : boolean;
  signal call_stmt_59_call_req_0 : boolean;
  signal call_stmt_59_call_ack_0 : boolean;
  signal call_stmt_59_call_req_1 : boolean;
  signal call_stmt_59_call_ack_1 : boolean;
  signal ADD_u8_u8_63_inst_req_0 : boolean;
  signal ADD_u8_u8_63_inst_ack_0 : boolean;
  signal ADD_u8_u8_63_inst_req_1 : boolean;
  signal ADD_u8_u8_63_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "add_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 80) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= rs1_data;
  rs1_data_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= rs2_data;
  rs2_data_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(71 downto 64) <= rd;
  rd_buffer <= in_buffer_data_out(71 downto 64);
  in_buffer_data_in(79 downto 72) <= pc;
  pc_buffer <= in_buffer_data_out(79 downto 72);
  in_buffer_data_in(tag_length + 79 downto 80) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 79 downto 80);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  add_CP_290_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "add_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= next_pc_buffer;
  next_pc <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= add_CP_290_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= add_CP_290_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= add_CP_290_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  add_CP_290: Block -- control-path 
    signal add_CP_290_elements: BooleanArray(7 downto 0);
    -- 
  begin -- 
    add_CP_290_elements(0) <= add_CP_290_start;
    add_CP_290_symbol <= add_CP_290_elements(7);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0:  members (17) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_54_to_assign_stmt_64/$entry
      -- CP-element group 0: 	 assign_stmt_54_to_assign_stmt_64/ADD_u32_u32_53_sample_start_
      -- CP-element group 0: 	 assign_stmt_54_to_assign_stmt_64/ADD_u32_u32_53_update_start_
      -- CP-element group 0: 	 assign_stmt_54_to_assign_stmt_64/ADD_u32_u32_53_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_54_to_assign_stmt_64/ADD_u32_u32_53_Sample/rr
      -- CP-element group 0: 	 assign_stmt_54_to_assign_stmt_64/ADD_u32_u32_53_Update/$entry
      -- CP-element group 0: 	 assign_stmt_54_to_assign_stmt_64/ADD_u32_u32_53_Update/cr
      -- CP-element group 0: 	 assign_stmt_54_to_assign_stmt_64/call_stmt_59_update_start_
      -- CP-element group 0: 	 assign_stmt_54_to_assign_stmt_64/call_stmt_59_Update/$entry
      -- CP-element group 0: 	 assign_stmt_54_to_assign_stmt_64/call_stmt_59_Update/ccr
      -- CP-element group 0: 	 assign_stmt_54_to_assign_stmt_64/ADD_u8_u8_63_sample_start_
      -- CP-element group 0: 	 assign_stmt_54_to_assign_stmt_64/ADD_u8_u8_63_update_start_
      -- CP-element group 0: 	 assign_stmt_54_to_assign_stmt_64/ADD_u8_u8_63_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_54_to_assign_stmt_64/ADD_u8_u8_63_Sample/rr
      -- CP-element group 0: 	 assign_stmt_54_to_assign_stmt_64/ADD_u8_u8_63_Update/$entry
      -- CP-element group 0: 	 assign_stmt_54_to_assign_stmt_64/ADD_u8_u8_63_Update/cr
      -- 
    rr_303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_CP_290_elements(0), ack => ADD_u32_u32_53_inst_req_0); -- 
    cr_308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_CP_290_elements(0), ack => ADD_u32_u32_53_inst_req_1); -- 
    ccr_322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_CP_290_elements(0), ack => call_stmt_59_call_req_1); -- 
    rr_331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_CP_290_elements(0), ack => ADD_u8_u8_63_inst_req_0); -- 
    cr_336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_CP_290_elements(0), ack => ADD_u8_u8_63_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_54_to_assign_stmt_64/ADD_u32_u32_53_sample_completed_
      -- CP-element group 1: 	 assign_stmt_54_to_assign_stmt_64/ADD_u32_u32_53_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_54_to_assign_stmt_64/ADD_u32_u32_53_Sample/ra
      -- 
    ra_304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_53_inst_ack_0, ack => add_CP_290_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_54_to_assign_stmt_64/ADD_u32_u32_53_update_completed_
      -- CP-element group 2: 	 assign_stmt_54_to_assign_stmt_64/ADD_u32_u32_53_Update/$exit
      -- CP-element group 2: 	 assign_stmt_54_to_assign_stmt_64/ADD_u32_u32_53_Update/ca
      -- CP-element group 2: 	 assign_stmt_54_to_assign_stmt_64/call_stmt_59_sample_start_
      -- CP-element group 2: 	 assign_stmt_54_to_assign_stmt_64/call_stmt_59_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_54_to_assign_stmt_64/call_stmt_59_Sample/crr
      -- 
    ca_309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_53_inst_ack_1, ack => add_CP_290_elements(2)); -- 
    crr_317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_CP_290_elements(2), ack => call_stmt_59_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_54_to_assign_stmt_64/call_stmt_59_sample_completed_
      -- CP-element group 3: 	 assign_stmt_54_to_assign_stmt_64/call_stmt_59_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_54_to_assign_stmt_64/call_stmt_59_Sample/cra
      -- 
    cra_318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_59_call_ack_0, ack => add_CP_290_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_54_to_assign_stmt_64/call_stmt_59_update_completed_
      -- CP-element group 4: 	 assign_stmt_54_to_assign_stmt_64/call_stmt_59_Update/$exit
      -- CP-element group 4: 	 assign_stmt_54_to_assign_stmt_64/call_stmt_59_Update/cca
      -- 
    cca_323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_59_call_ack_1, ack => add_CP_290_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_54_to_assign_stmt_64/ADD_u8_u8_63_sample_completed_
      -- CP-element group 5: 	 assign_stmt_54_to_assign_stmt_64/ADD_u8_u8_63_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_54_to_assign_stmt_64/ADD_u8_u8_63_Sample/ra
      -- 
    ra_332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_63_inst_ack_0, ack => add_CP_290_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_54_to_assign_stmt_64/ADD_u8_u8_63_update_completed_
      -- CP-element group 6: 	 assign_stmt_54_to_assign_stmt_64/ADD_u8_u8_63_Update/$exit
      -- CP-element group 6: 	 assign_stmt_54_to_assign_stmt_64/ADD_u8_u8_63_Update/ca
      -- 
    ca_337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_63_inst_ack_1, ack => add_CP_290_elements(6)); -- 
    -- CP-element group 7:  join  transition  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 $exit
      -- CP-element group 7: 	 assign_stmt_54_to_assign_stmt_64/$exit
      -- 
    add_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 22) := "add_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= add_CP_290_elements(4) & add_CP_290_elements(6);
      gj_add_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => add_CP_290_elements(7), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal dummy_59 : std_logic_vector(31 downto 0);
    signal konst_55_wire_constant : std_logic_vector(0 downto 0);
    signal konst_62_wire_constant : std_logic_vector(7 downto 0);
    signal output_54 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_55_wire_constant <= "0";
    konst_62_wire_constant <= "00000001";
    -- shared split operator group (0) : ADD_u32_u32_53_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= rs1_data_buffer & rs2_data_buffer;
      output_54 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_53_inst_req_0;
      ADD_u32_u32_53_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_53_inst_req_1;
      ADD_u32_u32_53_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : ADD_u8_u8_63_inst 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pc_buffer;
      next_pc_buffer <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_63_inst_req_0;
      ADD_u8_u8_63_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_63_inst_req_1;
      ADD_u8_u8_63_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared call operator group (0) : call_stmt_59_call 
    accessreg_call_group_0: Block -- 
      signal data_in: std_logic_vector(40 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_59_call_req_0;
      call_stmt_59_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_59_call_req_1;
      call_stmt_59_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessreg_call_group_0_gI: SplitGuardInterface generic map(name => "accessreg_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_55_wire_constant & rd_buffer & output_54;
      dummy_59 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 41,
        owidth => 41,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessreg_call_reqs(0),
          ackR => accessreg_call_acks(0),
          dataR => accessreg_call_data(40 downto 0),
          tagR => accessreg_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessreg_return_acks(0), -- cross-over
          ackL => accessreg_return_reqs(0), -- cross-over
          dataL => accessreg_return_data(31 downto 0),
          tagL => accessreg_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end add_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity and_i is -- 
  generic (tag_length : integer); 
  port ( -- 
    rs1_data : in  std_logic_vector(31 downto 0);
    rs2_data : in  std_logic_vector(31 downto 0);
    rd : in  std_logic_vector(7 downto 0);
    pc : in  std_logic_vector(7 downto 0);
    next_pc : out  std_logic_vector(7 downto 0);
    accessreg_call_reqs : out  std_logic_vector(0 downto 0);
    accessreg_call_acks : in   std_logic_vector(0 downto 0);
    accessreg_call_data : out  std_logic_vector(40 downto 0);
    accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
    accessreg_return_reqs : out  std_logic_vector(0 downto 0);
    accessreg_return_acks : in   std_logic_vector(0 downto 0);
    accessreg_return_data : in   std_logic_vector(31 downto 0);
    accessreg_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity and_i;
architecture and_i_arch of and_i is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 80)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rs1_data_buffer :  std_logic_vector(31 downto 0);
  signal rs1_data_update_enable: Boolean;
  signal rs2_data_buffer :  std_logic_vector(31 downto 0);
  signal rs2_data_update_enable: Boolean;
  signal rd_buffer :  std_logic_vector(7 downto 0);
  signal rd_update_enable: Boolean;
  signal pc_buffer :  std_logic_vector(7 downto 0);
  signal pc_update_enable: Boolean;
  -- output port buffer signals
  signal next_pc_buffer :  std_logic_vector(7 downto 0);
  signal next_pc_update_enable: Boolean;
  signal and_i_CP_338_start: Boolean;
  signal and_i_CP_338_symbol: Boolean;
  -- volatile/operator module components. 
  component accessreg is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(7 downto 0);
      write_data : in  std_logic_vector(31 downto 0);
      read_data : out  std_logic_vector(31 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal AND_u32_u32_75_inst_req_0 : boolean;
  signal AND_u32_u32_75_inst_ack_0 : boolean;
  signal AND_u32_u32_75_inst_req_1 : boolean;
  signal AND_u32_u32_75_inst_ack_1 : boolean;
  signal call_stmt_81_call_req_0 : boolean;
  signal call_stmt_81_call_ack_0 : boolean;
  signal call_stmt_81_call_req_1 : boolean;
  signal call_stmt_81_call_ack_1 : boolean;
  signal ADD_u8_u8_85_inst_req_0 : boolean;
  signal ADD_u8_u8_85_inst_ack_0 : boolean;
  signal ADD_u8_u8_85_inst_req_1 : boolean;
  signal ADD_u8_u8_85_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "and_i_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 80) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= rs1_data;
  rs1_data_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= rs2_data;
  rs2_data_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(71 downto 64) <= rd;
  rd_buffer <= in_buffer_data_out(71 downto 64);
  in_buffer_data_in(79 downto 72) <= pc;
  pc_buffer <= in_buffer_data_out(79 downto 72);
  in_buffer_data_in(tag_length + 79 downto 80) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 79 downto 80);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  and_i_CP_338_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "and_i_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= next_pc_buffer;
  next_pc <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= and_i_CP_338_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= and_i_CP_338_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= and_i_CP_338_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  and_i_CP_338: Block -- control-path 
    signal and_i_CP_338_elements: BooleanArray(7 downto 0);
    -- 
  begin -- 
    and_i_CP_338_elements(0) <= and_i_CP_338_start;
    and_i_CP_338_symbol <= and_i_CP_338_elements(7);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0:  members (17) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_76_to_assign_stmt_86/$entry
      -- CP-element group 0: 	 assign_stmt_76_to_assign_stmt_86/AND_u32_u32_75_sample_start_
      -- CP-element group 0: 	 assign_stmt_76_to_assign_stmt_86/AND_u32_u32_75_update_start_
      -- CP-element group 0: 	 assign_stmt_76_to_assign_stmt_86/AND_u32_u32_75_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_76_to_assign_stmt_86/AND_u32_u32_75_Sample/rr
      -- CP-element group 0: 	 assign_stmt_76_to_assign_stmt_86/AND_u32_u32_75_Update/$entry
      -- CP-element group 0: 	 assign_stmt_76_to_assign_stmt_86/AND_u32_u32_75_Update/cr
      -- CP-element group 0: 	 assign_stmt_76_to_assign_stmt_86/call_stmt_81_update_start_
      -- CP-element group 0: 	 assign_stmt_76_to_assign_stmt_86/call_stmt_81_Update/$entry
      -- CP-element group 0: 	 assign_stmt_76_to_assign_stmt_86/call_stmt_81_Update/ccr
      -- CP-element group 0: 	 assign_stmt_76_to_assign_stmt_86/ADD_u8_u8_85_sample_start_
      -- CP-element group 0: 	 assign_stmt_76_to_assign_stmt_86/ADD_u8_u8_85_update_start_
      -- CP-element group 0: 	 assign_stmt_76_to_assign_stmt_86/ADD_u8_u8_85_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_76_to_assign_stmt_86/ADD_u8_u8_85_Sample/rr
      -- CP-element group 0: 	 assign_stmt_76_to_assign_stmt_86/ADD_u8_u8_85_Update/$entry
      -- CP-element group 0: 	 assign_stmt_76_to_assign_stmt_86/ADD_u8_u8_85_Update/cr
      -- 
    rr_351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => and_i_CP_338_elements(0), ack => AND_u32_u32_75_inst_req_0); -- 
    cr_356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => and_i_CP_338_elements(0), ack => AND_u32_u32_75_inst_req_1); -- 
    ccr_370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => and_i_CP_338_elements(0), ack => call_stmt_81_call_req_1); -- 
    rr_379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => and_i_CP_338_elements(0), ack => ADD_u8_u8_85_inst_req_0); -- 
    cr_384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => and_i_CP_338_elements(0), ack => ADD_u8_u8_85_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_76_to_assign_stmt_86/AND_u32_u32_75_sample_completed_
      -- CP-element group 1: 	 assign_stmt_76_to_assign_stmt_86/AND_u32_u32_75_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_76_to_assign_stmt_86/AND_u32_u32_75_Sample/ra
      -- 
    ra_352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_75_inst_ack_0, ack => and_i_CP_338_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_76_to_assign_stmt_86/AND_u32_u32_75_update_completed_
      -- CP-element group 2: 	 assign_stmt_76_to_assign_stmt_86/AND_u32_u32_75_Update/$exit
      -- CP-element group 2: 	 assign_stmt_76_to_assign_stmt_86/AND_u32_u32_75_Update/ca
      -- CP-element group 2: 	 assign_stmt_76_to_assign_stmt_86/call_stmt_81_sample_start_
      -- CP-element group 2: 	 assign_stmt_76_to_assign_stmt_86/call_stmt_81_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_76_to_assign_stmt_86/call_stmt_81_Sample/crr
      -- 
    ca_357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_75_inst_ack_1, ack => and_i_CP_338_elements(2)); -- 
    crr_365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => and_i_CP_338_elements(2), ack => call_stmt_81_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_76_to_assign_stmt_86/call_stmt_81_sample_completed_
      -- CP-element group 3: 	 assign_stmt_76_to_assign_stmt_86/call_stmt_81_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_76_to_assign_stmt_86/call_stmt_81_Sample/cra
      -- 
    cra_366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_81_call_ack_0, ack => and_i_CP_338_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_76_to_assign_stmt_86/call_stmt_81_update_completed_
      -- CP-element group 4: 	 assign_stmt_76_to_assign_stmt_86/call_stmt_81_Update/$exit
      -- CP-element group 4: 	 assign_stmt_76_to_assign_stmt_86/call_stmt_81_Update/cca
      -- 
    cca_371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_81_call_ack_1, ack => and_i_CP_338_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_76_to_assign_stmt_86/ADD_u8_u8_85_sample_completed_
      -- CP-element group 5: 	 assign_stmt_76_to_assign_stmt_86/ADD_u8_u8_85_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_76_to_assign_stmt_86/ADD_u8_u8_85_Sample/ra
      -- 
    ra_380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_85_inst_ack_0, ack => and_i_CP_338_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_76_to_assign_stmt_86/ADD_u8_u8_85_update_completed_
      -- CP-element group 6: 	 assign_stmt_76_to_assign_stmt_86/ADD_u8_u8_85_Update/$exit
      -- CP-element group 6: 	 assign_stmt_76_to_assign_stmt_86/ADD_u8_u8_85_Update/ca
      -- 
    ca_385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_85_inst_ack_1, ack => and_i_CP_338_elements(6)); -- 
    -- CP-element group 7:  join  transition  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 $exit
      -- CP-element group 7: 	 assign_stmt_76_to_assign_stmt_86/$exit
      -- 
    and_i_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "and_i_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= and_i_CP_338_elements(4) & and_i_CP_338_elements(6);
      gj_and_i_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => and_i_CP_338_elements(7), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal dummy1_81 : std_logic_vector(31 downto 0);
    signal konst_77_wire_constant : std_logic_vector(0 downto 0);
    signal konst_84_wire_constant : std_logic_vector(7 downto 0);
    signal output_76 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_77_wire_constant <= "0";
    konst_84_wire_constant <= "00000001";
    -- shared split operator group (0) : ADD_u8_u8_85_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pc_buffer;
      next_pc_buffer <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_85_inst_req_0;
      ADD_u8_u8_85_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_85_inst_req_1;
      ADD_u8_u8_85_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : AND_u32_u32_75_inst 
    ApIntAnd_group_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= rs1_data_buffer & rs2_data_buffer;
      output_76 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_75_inst_req_0;
      AND_u32_u32_75_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_75_inst_req_1;
      AND_u32_u32_75_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared call operator group (0) : call_stmt_81_call 
    accessreg_call_group_0: Block -- 
      signal data_in: std_logic_vector(40 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_81_call_req_0;
      call_stmt_81_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_81_call_req_1;
      call_stmt_81_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessreg_call_group_0_gI: SplitGuardInterface generic map(name => "accessreg_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_77_wire_constant & rd_buffer & output_76;
      dummy1_81 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 41,
        owidth => 41,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessreg_call_reqs(0),
          ackR => accessreg_call_acks(0),
          dataR => accessreg_call_data(40 downto 0),
          tagR => accessreg_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessreg_return_acks(0), -- cross-over
          ackL => accessreg_return_reqs(0), -- cross-over
          dataL => accessreg_return_data(31 downto 0),
          tagL => accessreg_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end and_i_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity bn is -- 
  generic (tag_length : integer); 
  port ( -- 
    rs1_data : in  std_logic_vector(31 downto 0);
    rs2_data : in  std_logic_vector(31 downto 0);
    rd : in  std_logic_vector(7 downto 0);
    pc : in  std_logic_vector(7 downto 0);
    next_pc : out  std_logic_vector(7 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity bn;
architecture bn_arch of bn is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 80)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rs1_data_buffer :  std_logic_vector(31 downto 0);
  signal rs1_data_update_enable: Boolean;
  signal rs2_data_buffer :  std_logic_vector(31 downto 0);
  signal rs2_data_update_enable: Boolean;
  signal rd_buffer :  std_logic_vector(7 downto 0);
  signal rd_update_enable: Boolean;
  signal pc_buffer :  std_logic_vector(7 downto 0);
  signal pc_update_enable: Boolean;
  -- output port buffer signals
  signal next_pc_buffer :  std_logic_vector(7 downto 0);
  signal next_pc_update_enable: Boolean;
  signal bn_CP_386_start: Boolean;
  signal bn_CP_386_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LSHR_u32_u32_97_inst_req_0 : boolean;
  signal LSHR_u32_u32_97_inst_ack_0 : boolean;
  signal LSHR_u32_u32_97_inst_req_1 : boolean;
  signal LSHR_u32_u32_97_inst_ack_1 : boolean;
  signal ADD_u8_u8_103_inst_req_0 : boolean;
  signal ADD_u8_u8_103_inst_ack_0 : boolean;
  signal ADD_u8_u8_103_inst_req_1 : boolean;
  signal ADD_u8_u8_103_inst_ack_1 : boolean;
  signal STORE_next_pc1_100_store_0_req_0 : boolean;
  signal STORE_next_pc1_100_store_0_ack_0 : boolean;
  signal STORE_next_pc1_100_store_0_req_1 : boolean;
  signal STORE_next_pc1_100_store_0_ack_1 : boolean;
  signal slice_108_inst_req_0 : boolean;
  signal slice_108_inst_ack_0 : boolean;
  signal slice_108_inst_req_1 : boolean;
  signal slice_108_inst_ack_1 : boolean;
  signal STORE_next_pc1_106_store_0_req_0 : boolean;
  signal STORE_next_pc1_106_store_0_ack_0 : boolean;
  signal STORE_next_pc1_106_store_0_req_1 : boolean;
  signal STORE_next_pc1_106_store_0_ack_1 : boolean;
  signal LOAD_next_pc1_111_load_0_req_0 : boolean;
  signal LOAD_next_pc1_111_load_0_ack_0 : boolean;
  signal LOAD_next_pc1_111_load_0_req_1 : boolean;
  signal LOAD_next_pc1_111_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "bn_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 80) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= rs1_data;
  rs1_data_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= rs2_data;
  rs2_data_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(71 downto 64) <= rd;
  rd_buffer <= in_buffer_data_out(71 downto 64);
  in_buffer_data_in(79 downto 72) <= pc;
  pc_buffer <= in_buffer_data_out(79 downto 72);
  in_buffer_data_in(tag_length + 79 downto 80) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 79 downto 80);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  bn_CP_386_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "bn_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= next_pc_buffer;
  next_pc <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= bn_CP_386_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= bn_CP_386_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= bn_CP_386_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  bn_CP_386: Block -- control-path 
    signal bn_CP_386_elements: BooleanArray(18 downto 0);
    -- 
  begin -- 
    bn_CP_386_elements(0) <= bn_CP_386_start;
    bn_CP_386_symbol <= bn_CP_386_elements(18);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	10 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	15 
    -- CP-element group 0:  members (35) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/$entry
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/LSHR_u32_u32_97_sample_start_
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/LSHR_u32_u32_97_update_start_
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/LSHR_u32_u32_97_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/LSHR_u32_u32_97_Sample/rr
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/LSHR_u32_u32_97_Update/$entry
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/LSHR_u32_u32_97_Update/cr
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/ADD_u8_u8_103_update_start_
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/ADD_u8_u8_103_Update/$entry
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/ADD_u8_u8_103_Update/cr
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_update_start_
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_Update/$entry
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/slice_108_update_start_
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/slice_108_Update/$entry
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/slice_108_Update/cr
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_update_start_
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_Update/$entry
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_update_start_
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_Update/$entry
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_Update/word_access_complete/word_0/cr
      -- 
    rr_399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bn_CP_386_elements(0), ack => LSHR_u32_u32_97_inst_req_0); -- 
    cr_404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bn_CP_386_elements(0), ack => LSHR_u32_u32_97_inst_req_1); -- 
    cr_418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bn_CP_386_elements(0), ack => ADD_u8_u8_103_inst_req_1); -- 
    cr_451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bn_CP_386_elements(0), ack => STORE_next_pc1_100_store_0_req_1); -- 
    cr_465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bn_CP_386_elements(0), ack => slice_108_inst_req_1); -- 
    cr_498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bn_CP_386_elements(0), ack => STORE_next_pc1_106_store_0_req_1); -- 
    cr_526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bn_CP_386_elements(0), ack => LOAD_next_pc1_111_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_98_to_assign_stmt_112/LSHR_u32_u32_97_sample_completed_
      -- CP-element group 1: 	 assign_stmt_98_to_assign_stmt_112/LSHR_u32_u32_97_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_98_to_assign_stmt_112/LSHR_u32_u32_97_Sample/ra
      -- 
    ra_400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_97_inst_ack_0, ack => bn_CP_386_elements(1)); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 assign_stmt_98_to_assign_stmt_112/LSHR_u32_u32_97_update_completed_
      -- CP-element group 2: 	 assign_stmt_98_to_assign_stmt_112/LSHR_u32_u32_97_Update/$exit
      -- CP-element group 2: 	 assign_stmt_98_to_assign_stmt_112/LSHR_u32_u32_97_Update/ca
      -- CP-element group 2: 	 assign_stmt_98_to_assign_stmt_112/ADD_u8_u8_103_sample_start_
      -- CP-element group 2: 	 assign_stmt_98_to_assign_stmt_112/ADD_u8_u8_103_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_98_to_assign_stmt_112/ADD_u8_u8_103_Sample/rr
      -- CP-element group 2: 	 assign_stmt_98_to_assign_stmt_112/slice_108_sample_start_
      -- CP-element group 2: 	 assign_stmt_98_to_assign_stmt_112/slice_108_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_98_to_assign_stmt_112/slice_108_Sample/rr
      -- 
    ca_405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_97_inst_ack_1, ack => bn_CP_386_elements(2)); -- 
    rr_413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bn_CP_386_elements(2), ack => ADD_u8_u8_103_inst_req_0); -- 
    rr_460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bn_CP_386_elements(2), ack => slice_108_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_98_to_assign_stmt_112/ADD_u8_u8_103_sample_completed_
      -- CP-element group 3: 	 assign_stmt_98_to_assign_stmt_112/ADD_u8_u8_103_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_98_to_assign_stmt_112/ADD_u8_u8_103_Sample/ra
      -- 
    ra_414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_103_inst_ack_0, ack => bn_CP_386_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_98_to_assign_stmt_112/ADD_u8_u8_103_update_completed_
      -- CP-element group 4: 	 assign_stmt_98_to_assign_stmt_112/ADD_u8_u8_103_Update/$exit
      -- CP-element group 4: 	 assign_stmt_98_to_assign_stmt_112/ADD_u8_u8_103_Update/ca
      -- 
    ca_419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_103_inst_ack_1, ack => bn_CP_386_elements(4)); -- 
    -- CP-element group 5:  join  transition  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (9) 
      -- CP-element group 5: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_sample_start_
      -- CP-element group 5: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_Sample/$entry
      -- CP-element group 5: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_Sample/STORE_next_pc1_100_Split/$entry
      -- CP-element group 5: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_Sample/STORE_next_pc1_100_Split/$exit
      -- CP-element group 5: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_Sample/STORE_next_pc1_100_Split/split_req
      -- CP-element group 5: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_Sample/STORE_next_pc1_100_Split/split_ack
      -- CP-element group 5: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_Sample/word_access_start/$entry
      -- CP-element group 5: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_Sample/word_access_start/word_0/$entry
      -- CP-element group 5: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_Sample/word_access_start/word_0/rr
      -- 
    rr_440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bn_CP_386_elements(5), ack => STORE_next_pc1_100_store_0_req_0); -- 
    bn_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 21) := "bn_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= bn_CP_386_elements(0) & bn_CP_386_elements(2) & bn_CP_386_elements(4);
      gj_bn_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => bn_CP_386_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	16 
    -- CP-element group 6:  members (5) 
      -- CP-element group 6: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_sample_completed_
      -- CP-element group 6: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_Sample/$exit
      -- CP-element group 6: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_Sample/word_access_start/$exit
      -- CP-element group 6: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_Sample/word_access_start/word_0/$exit
      -- CP-element group 6: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_Sample/word_access_start/word_0/ra
      -- 
    ra_441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_next_pc1_100_store_0_ack_0, ack => bn_CP_386_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	18 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_update_completed_
      -- CP-element group 7: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_Update/$exit
      -- CP-element group 7: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_Update/word_access_complete/$exit
      -- CP-element group 7: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_Update/word_access_complete/word_0/$exit
      -- CP-element group 7: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_Update/word_access_complete/word_0/ca
      -- 
    ca_452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_next_pc1_100_store_0_ack_1, ack => bn_CP_386_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_98_to_assign_stmt_112/slice_108_sample_completed_
      -- CP-element group 8: 	 assign_stmt_98_to_assign_stmt_112/slice_108_Sample/$exit
      -- CP-element group 8: 	 assign_stmt_98_to_assign_stmt_112/slice_108_Sample/ra
      -- 
    ra_461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_108_inst_ack_0, ack => bn_CP_386_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_98_to_assign_stmt_112/slice_108_update_completed_
      -- CP-element group 9: 	 assign_stmt_98_to_assign_stmt_112/slice_108_Update/$exit
      -- CP-element group 9: 	 assign_stmt_98_to_assign_stmt_112/slice_108_Update/ca
      -- 
    ca_466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_108_inst_ack_1, ack => bn_CP_386_elements(9)); -- 
    -- CP-element group 10:  join  transition  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: 	9 
    -- CP-element group 10: 	16 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_sample_start_
      -- CP-element group 10: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_Sample/STORE_next_pc1_106_Split/$entry
      -- CP-element group 10: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_Sample/STORE_next_pc1_106_Split/$exit
      -- CP-element group 10: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_Sample/STORE_next_pc1_106_Split/split_req
      -- CP-element group 10: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_Sample/STORE_next_pc1_106_Split/split_ack
      -- CP-element group 10: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_Sample/word_access_start/$entry
      -- CP-element group 10: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_Sample/word_access_start/word_0/$entry
      -- CP-element group 10: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_Sample/word_access_start/word_0/rr
      -- 
    rr_487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bn_CP_386_elements(10), ack => STORE_next_pc1_106_store_0_req_0); -- 
    bn_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 22) := "bn_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= bn_CP_386_elements(0) & bn_CP_386_elements(9) & bn_CP_386_elements(16);
      gj_bn_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => bn_CP_386_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_sample_completed_
      -- CP-element group 11: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_Sample/$exit
      -- CP-element group 11: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_Sample/word_access_start/$exit
      -- CP-element group 11: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_Sample/word_access_start/word_0/ra
      -- 
    ra_488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_next_pc1_106_store_0_ack_0, ack => bn_CP_386_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	18 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_update_completed_
      -- CP-element group 12: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_Update/$exit
      -- CP-element group 12: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_Update/word_access_complete/$exit
      -- CP-element group 12: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_Update/word_access_complete/word_0/ca
      -- 
    ca_499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_next_pc1_106_store_0_ack_1, ack => bn_CP_386_elements(12)); -- 
    -- CP-element group 13:  join  transition  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: 	17 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_sample_start_
      -- CP-element group 13: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_Sample/$entry
      -- CP-element group 13: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_Sample/word_access_start/$entry
      -- CP-element group 13: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_Sample/word_access_start/word_0/$entry
      -- CP-element group 13: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_Sample/word_access_start/word_0/rr
      -- 
    rr_515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bn_CP_386_elements(13), ack => LOAD_next_pc1_111_load_0_req_0); -- 
    bn_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 22) := "bn_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= bn_CP_386_elements(0) & bn_CP_386_elements(17);
      gj_bn_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => bn_CP_386_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (5) 
      -- CP-element group 14: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_sample_completed_
      -- CP-element group 14: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_Sample/$exit
      -- CP-element group 14: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_Sample/word_access_start/$exit
      -- CP-element group 14: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_Sample/word_access_start/word_0/$exit
      -- CP-element group 14: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_Sample/word_access_start/word_0/ra
      -- 
    ra_516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_next_pc1_111_load_0_ack_0, ack => bn_CP_386_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	0 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	18 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_update_completed_
      -- CP-element group 15: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_Update/$exit
      -- CP-element group 15: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_Update/word_access_complete/$exit
      -- CP-element group 15: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_Update/word_access_complete/word_0/$exit
      -- CP-element group 15: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_Update/word_access_complete/word_0/ca
      -- CP-element group 15: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_Update/LOAD_next_pc1_111_Merge/$entry
      -- CP-element group 15: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_Update/LOAD_next_pc1_111_Merge/$exit
      -- CP-element group 15: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_Update/LOAD_next_pc1_111_Merge/merge_req
      -- CP-element group 15: 	 assign_stmt_98_to_assign_stmt_112/LOAD_next_pc1_111_Update/LOAD_next_pc1_111_Merge/merge_ack
      -- 
    ca_527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_next_pc1_111_load_0_ack_1, ack => bn_CP_386_elements(15)); -- 
    -- CP-element group 16:  transition  delay-element  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	6 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	10 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_100_STORE_next_pc1_106_delay
      -- 
    -- Element group bn_CP_386_elements(16) is a control-delay.
    cp_element_16_delay: control_delay_element  generic map(name => " 16_delay", delay_value => 1)  port map(req => bn_CP_386_elements(6), ack => bn_CP_386_elements(16), clk => clk, reset =>reset);
    -- CP-element group 17:  transition  delay-element  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	13 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 assign_stmt_98_to_assign_stmt_112/STORE_next_pc1_106_LOAD_next_pc1_111_delay
      -- 
    -- Element group bn_CP_386_elements(17) is a control-delay.
    cp_element_17_delay: control_delay_element  generic map(name => " 17_delay", delay_value => 1)  port map(req => bn_CP_386_elements(11), ack => bn_CP_386_elements(17), clk => clk, reset =>reset);
    -- CP-element group 18:  join  transition  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	7 
    -- CP-element group 18: 	12 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 $exit
      -- CP-element group 18: 	 assign_stmt_98_to_assign_stmt_112/$exit
      -- 
    bn_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 22) := "bn_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= bn_CP_386_elements(7) & bn_CP_386_elements(12) & bn_CP_386_elements(15);
      gj_bn_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => bn_CP_386_elements(18), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u8_u8_103_wire : std_logic_vector(7 downto 0);
    signal LOAD_next_pc1_111_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_next_pc1_111_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_next_pc1_100_data_0 : std_logic_vector(7 downto 0);
    signal STORE_next_pc1_100_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_next_pc1_106_data_0 : std_logic_vector(7 downto 0);
    signal STORE_next_pc1_106_word_address_0 : std_logic_vector(0 downto 0);
    signal bnn_98 : std_logic_vector(31 downto 0);
    signal konst_102_wire_constant : std_logic_vector(7 downto 0);
    signal konst_96_wire_constant : std_logic_vector(31 downto 0);
    signal slice_108_wire : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    LOAD_next_pc1_111_word_address_0 <= "0";
    STORE_next_pc1_100_word_address_0 <= "0";
    STORE_next_pc1_106_word_address_0 <= "0";
    konst_102_wire_constant <= "00000001";
    konst_96_wire_constant <= "00000000000000000000000000011111";
    slice_108_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      signal sample_req_ug, sample_ack_ug, update_req_ug, update_ack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      sample_req_ug(0) <= slice_108_inst_req_0;
      slice_108_inst_ack_0<= sample_ack_ug(0);
      update_req_ug(0) <= slice_108_inst_req_1;
      slice_108_inst_ack_1<= update_ack_ug(0);
      guard_vector(0) <=  bnn_98(0);
      slice_108_inst_gI: SplitGuardInterface generic map(name => "slice_108_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_ug,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_ug,
        cr_in => update_req_ug,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_ug,
        guards => guard_vector); -- 
      slice_108_inst: SliceSplitProtocol generic map(name => "slice_108_inst", in_data_width => 32, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => rs2_data_buffer, dout => slice_108_wire, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- equivalence LOAD_next_pc1_111_gather_scatter
    process(LOAD_next_pc1_111_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_next_pc1_111_data_0;
      ov(7 downto 0) := iv;
      next_pc_buffer <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_next_pc1_100_gather_scatter
    process(ADD_u8_u8_103_wire) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u8_u8_103_wire;
      ov(7 downto 0) := iv;
      STORE_next_pc1_100_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_next_pc1_106_gather_scatter
    process(slice_108_wire) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := slice_108_wire;
      ov(7 downto 0) := iv;
      STORE_next_pc1_106_data_0 <= ov(7 downto 0);
      --
    end process;
    -- shared split operator group (0) : ADD_u8_u8_103_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pc_buffer;
      ADD_u8_u8_103_wire <= data_out(7 downto 0);
      guard_vector(0)  <=  not bnn_98(0);
      reqL_unguarded(0) <= ADD_u8_u8_103_inst_req_0;
      ADD_u8_u8_103_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_103_inst_req_1;
      ADD_u8_u8_103_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : LSHR_u32_u32_97_inst 
    ApIntLSHR_group_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= rs1_data_buffer;
      bnn_98 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_97_inst_req_0;
      LSHR_u32_u32_97_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_97_inst_req_1;
      LSHR_u32_u32_97_inst_ack_1 <= ackR_unguarded(0);
      ApIntLSHR_group_1_gI: SplitGuardInterface generic map(name => "ApIntLSHR_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000011111",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared load operator group (0) : LOAD_next_pc1_111_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_next_pc1_111_load_0_req_0;
      LOAD_next_pc1_111_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_next_pc1_111_load_0_req_1;
      LOAD_next_pc1_111_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_next_pc1_111_word_address_0;
      LOAD_next_pc1_111_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(0 downto 0),
          mtag => memory_space_1_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(7 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : STORE_next_pc1_100_store_0 STORE_next_pc1_106_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(1 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= STORE_next_pc1_100_store_0_req_0;
      reqL_unguarded(0) <= STORE_next_pc1_106_store_0_req_0;
      STORE_next_pc1_100_store_0_ack_0 <= ackL_unguarded(1);
      STORE_next_pc1_106_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= STORE_next_pc1_100_store_0_req_1;
      reqR_unguarded(0) <= STORE_next_pc1_106_store_0_req_1;
      STORE_next_pc1_100_store_0_ack_1 <= ackR_unguarded(1);
      STORE_next_pc1_106_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= bnn_98(0);
      guard_vector(1)  <=  not bnn_98(0);
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_next_pc1_100_word_address_0 & STORE_next_pc1_106_word_address_0;
      data_in <= STORE_next_pc1_100_data_0 & STORE_next_pc1_106_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(0 downto 0),
          mdata => memory_space_1_sr_data(7 downto 0),
          mtag => memory_space_1_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end bn_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity bz is -- 
  generic (tag_length : integer); 
  port ( -- 
    rs1_data : in  std_logic_vector(31 downto 0);
    rs2_data : in  std_logic_vector(31 downto 0);
    rd : in  std_logic_vector(7 downto 0);
    pc : in  std_logic_vector(7 downto 0);
    next_pc : out  std_logic_vector(7 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity bz;
architecture bz_arch of bz is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 80)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rs1_data_buffer :  std_logic_vector(31 downto 0);
  signal rs1_data_update_enable: Boolean;
  signal rs2_data_buffer :  std_logic_vector(31 downto 0);
  signal rs2_data_update_enable: Boolean;
  signal rd_buffer :  std_logic_vector(7 downto 0);
  signal rd_update_enable: Boolean;
  signal pc_buffer :  std_logic_vector(7 downto 0);
  signal pc_update_enable: Boolean;
  -- output port buffer signals
  signal next_pc_buffer :  std_logic_vector(7 downto 0);
  signal next_pc_update_enable: Boolean;
  signal bz_CP_535_start: Boolean;
  signal bz_CP_535_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal W_bzz_120_inst_ack_1 : boolean;
  signal LOAD_next_pc1_135_load_0_ack_1 : boolean;
  signal LOAD_next_pc1_135_load_0_req_1 : boolean;
  signal W_bzz_120_inst_req_1 : boolean;
  signal STORE_next_pc1_124_store_0_ack_1 : boolean;
  signal STORE_next_pc1_124_store_0_req_1 : boolean;
  signal W_bzz_120_inst_ack_0 : boolean;
  signal LOAD_next_pc1_135_load_0_ack_0 : boolean;
  signal LOAD_next_pc1_135_load_0_req_0 : boolean;
  signal STORE_next_pc1_130_store_0_ack_1 : boolean;
  signal STORE_next_pc1_130_store_0_req_1 : boolean;
  signal ADD_u8_u8_127_inst_ack_1 : boolean;
  signal ADD_u8_u8_127_inst_req_1 : boolean;
  signal STORE_next_pc1_124_store_0_ack_0 : boolean;
  signal ADD_u8_u8_127_inst_ack_0 : boolean;
  signal STORE_next_pc1_124_store_0_req_0 : boolean;
  signal ADD_u8_u8_127_inst_req_0 : boolean;
  signal W_bzz_120_inst_req_0 : boolean;
  signal STORE_next_pc1_130_store_0_ack_0 : boolean;
  signal STORE_next_pc1_130_store_0_req_0 : boolean;
  signal slice_132_inst_ack_1 : boolean;
  signal slice_132_inst_req_1 : boolean;
  signal slice_132_inst_ack_0 : boolean;
  signal slice_132_inst_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "bz_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 80) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= rs1_data;
  rs1_data_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= rs2_data;
  rs2_data_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(71 downto 64) <= rd;
  rd_buffer <= in_buffer_data_out(71 downto 64);
  in_buffer_data_in(79 downto 72) <= pc;
  pc_buffer <= in_buffer_data_out(79 downto 72);
  in_buffer_data_in(tag_length + 79 downto 80) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 79 downto 80);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  bz_CP_535_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "bz_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= next_pc_buffer;
  next_pc <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= bz_CP_535_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= bz_CP_535_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= bz_CP_535_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  bz_CP_535: Block -- control-path 
    signal bz_CP_535_elements: BooleanArray(18 downto 0);
    -- 
  begin -- 
    bz_CP_535_elements(0) <= bz_CP_535_start;
    bz_CP_535_symbol <= bz_CP_535_elements(18);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	10 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	15 
    -- CP-element group 0:  members (35) 
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/$entry
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/assign_stmt_122_Update/req
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/assign_stmt_122_Update/$entry
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_Update/$entry
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/assign_stmt_122_update_start_
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/assign_stmt_122_sample_start_
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/ADD_u8_u8_127_update_start_
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_update_start_
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_update_start_
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_update_start_
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/ADD_u8_u8_127_Update/cr
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_Update/$entry
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/ADD_u8_u8_127_Update/$entry
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_Update/$entry
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/assign_stmt_122_Sample/req
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/assign_stmt_122_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/slice_132_Update/cr
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/slice_132_Update/$entry
      -- CP-element group 0: 	 assign_stmt_122_to_assign_stmt_136/slice_132_update_start_
      -- 
    req_548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bz_CP_535_elements(0), ack => W_bzz_120_inst_req_0); -- 
    req_553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bz_CP_535_elements(0), ack => W_bzz_120_inst_req_1); -- 
    cr_567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bz_CP_535_elements(0), ack => ADD_u8_u8_127_inst_req_1); -- 
    cr_600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bz_CP_535_elements(0), ack => STORE_next_pc1_124_store_0_req_1); -- 
    cr_614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bz_CP_535_elements(0), ack => slice_132_inst_req_1); -- 
    cr_647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bz_CP_535_elements(0), ack => STORE_next_pc1_130_store_0_req_1); -- 
    cr_675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bz_CP_535_elements(0), ack => LOAD_next_pc1_135_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_122_to_assign_stmt_136/assign_stmt_122_Sample/ack
      -- CP-element group 1: 	 assign_stmt_122_to_assign_stmt_136/assign_stmt_122_sample_completed_
      -- CP-element group 1: 	 assign_stmt_122_to_assign_stmt_136/assign_stmt_122_Sample/$exit
      -- 
    ack_549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bzz_120_inst_ack_0, ack => bz_CP_535_elements(1)); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 assign_stmt_122_to_assign_stmt_136/assign_stmt_122_Update/ack
      -- CP-element group 2: 	 assign_stmt_122_to_assign_stmt_136/ADD_u8_u8_127_sample_start_
      -- CP-element group 2: 	 assign_stmt_122_to_assign_stmt_136/ADD_u8_u8_127_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_122_to_assign_stmt_136/slice_132_sample_start_
      -- CP-element group 2: 	 assign_stmt_122_to_assign_stmt_136/assign_stmt_122_Update/$exit
      -- CP-element group 2: 	 assign_stmt_122_to_assign_stmt_136/ADD_u8_u8_127_Sample/rr
      -- CP-element group 2: 	 assign_stmt_122_to_assign_stmt_136/assign_stmt_122_update_completed_
      -- CP-element group 2: 	 assign_stmt_122_to_assign_stmt_136/slice_132_Sample/rr
      -- CP-element group 2: 	 assign_stmt_122_to_assign_stmt_136/slice_132_Sample/$entry
      -- 
    ack_554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bzz_120_inst_ack_1, ack => bz_CP_535_elements(2)); -- 
    rr_562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bz_CP_535_elements(2), ack => ADD_u8_u8_127_inst_req_0); -- 
    rr_609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bz_CP_535_elements(2), ack => slice_132_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_122_to_assign_stmt_136/ADD_u8_u8_127_sample_completed_
      -- CP-element group 3: 	 assign_stmt_122_to_assign_stmt_136/ADD_u8_u8_127_Sample/ra
      -- CP-element group 3: 	 assign_stmt_122_to_assign_stmt_136/ADD_u8_u8_127_Sample/$exit
      -- 
    ra_563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_127_inst_ack_0, ack => bz_CP_535_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_122_to_assign_stmt_136/ADD_u8_u8_127_update_completed_
      -- CP-element group 4: 	 assign_stmt_122_to_assign_stmt_136/ADD_u8_u8_127_Update/ca
      -- CP-element group 4: 	 assign_stmt_122_to_assign_stmt_136/ADD_u8_u8_127_Update/$exit
      -- 
    ca_568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_127_inst_ack_1, ack => bz_CP_535_elements(4)); -- 
    -- CP-element group 5:  join  transition  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (9) 
      -- CP-element group 5: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_Sample/word_access_start/$entry
      -- CP-element group 5: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_Sample/STORE_next_pc1_124_Split/split_ack
      -- CP-element group 5: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_Sample/STORE_next_pc1_124_Split/split_req
      -- CP-element group 5: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_Sample/STORE_next_pc1_124_Split/$exit
      -- CP-element group 5: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_Sample/STORE_next_pc1_124_Split/$entry
      -- CP-element group 5: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_Sample/$entry
      -- CP-element group 5: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_sample_start_
      -- CP-element group 5: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_Sample/word_access_start/word_0/rr
      -- CP-element group 5: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_Sample/word_access_start/word_0/$entry
      -- 
    rr_589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bz_CP_535_elements(5), ack => STORE_next_pc1_124_store_0_req_0); -- 
    bz_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 21) := "bz_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= bz_CP_535_elements(0) & bz_CP_535_elements(2) & bz_CP_535_elements(4);
      gj_bz_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => bz_CP_535_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	16 
    -- CP-element group 6:  members (5) 
      -- CP-element group 6: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_Sample/word_access_start/$exit
      -- CP-element group 6: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_Sample/$exit
      -- CP-element group 6: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_sample_completed_
      -- CP-element group 6: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_Sample/word_access_start/word_0/ra
      -- CP-element group 6: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_Sample/word_access_start/word_0/$exit
      -- 
    ra_590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_next_pc1_124_store_0_ack_0, ack => bz_CP_535_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	18 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_Update/word_access_complete/word_0/ca
      -- CP-element group 7: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_Update/word_access_complete/word_0/$exit
      -- CP-element group 7: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_Update/word_access_complete/$exit
      -- CP-element group 7: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_update_completed_
      -- CP-element group 7: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_Update/$exit
      -- 
    ca_601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_next_pc1_124_store_0_ack_1, ack => bz_CP_535_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_122_to_assign_stmt_136/slice_132_Sample/ra
      -- CP-element group 8: 	 assign_stmt_122_to_assign_stmt_136/slice_132_Sample/$exit
      -- CP-element group 8: 	 assign_stmt_122_to_assign_stmt_136/slice_132_sample_completed_
      -- 
    ra_610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_132_inst_ack_0, ack => bz_CP_535_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_122_to_assign_stmt_136/slice_132_Update/ca
      -- CP-element group 9: 	 assign_stmt_122_to_assign_stmt_136/slice_132_Update/$exit
      -- CP-element group 9: 	 assign_stmt_122_to_assign_stmt_136/slice_132_update_completed_
      -- 
    ca_615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_132_inst_ack_1, ack => bz_CP_535_elements(9)); -- 
    -- CP-element group 10:  join  transition  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: 	9 
    -- CP-element group 10: 	16 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_sample_start_
      -- CP-element group 10: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_Sample/word_access_start/word_0/rr
      -- CP-element group 10: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_Sample/word_access_start/word_0/$entry
      -- CP-element group 10: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_Sample/word_access_start/$entry
      -- CP-element group 10: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_Sample/STORE_next_pc1_130_Split/split_ack
      -- CP-element group 10: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_Sample/STORE_next_pc1_130_Split/split_req
      -- CP-element group 10: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_Sample/STORE_next_pc1_130_Split/$exit
      -- CP-element group 10: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_Sample/STORE_next_pc1_130_Split/$entry
      -- CP-element group 10: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_Sample/$entry
      -- 
    rr_636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bz_CP_535_elements(10), ack => STORE_next_pc1_130_store_0_req_0); -- 
    bz_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 22) := "bz_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= bz_CP_535_elements(0) & bz_CP_535_elements(9) & bz_CP_535_elements(16);
      gj_bz_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => bz_CP_535_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_sample_completed_
      -- CP-element group 11: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_Sample/word_access_start/word_0/ra
      -- CP-element group 11: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_Sample/word_access_start/$exit
      -- CP-element group 11: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_Sample/$exit
      -- 
    ra_637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_next_pc1_130_store_0_ack_0, ack => bz_CP_535_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	18 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_Update/word_access_complete/$exit
      -- CP-element group 12: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_Update/$exit
      -- CP-element group 12: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_update_completed_
      -- 
    ca_648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_next_pc1_130_store_0_ack_1, ack => bz_CP_535_elements(12)); -- 
    -- CP-element group 13:  join  transition  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: 	17 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_Sample/word_access_start/word_0/rr
      -- CP-element group 13: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_Sample/word_access_start/word_0/$entry
      -- CP-element group 13: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_Sample/word_access_start/$entry
      -- CP-element group 13: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_Sample/$entry
      -- CP-element group 13: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_sample_start_
      -- 
    rr_664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => bz_CP_535_elements(13), ack => LOAD_next_pc1_135_load_0_req_0); -- 
    bz_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 22) := "bz_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= bz_CP_535_elements(0) & bz_CP_535_elements(17);
      gj_bz_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => bz_CP_535_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (5) 
      -- CP-element group 14: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_Sample/word_access_start/word_0/ra
      -- CP-element group 14: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_Sample/word_access_start/word_0/$exit
      -- CP-element group 14: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_Sample/word_access_start/$exit
      -- CP-element group 14: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_Sample/$exit
      -- CP-element group 14: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_sample_completed_
      -- 
    ra_665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_next_pc1_135_load_0_ack_0, ack => bz_CP_535_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	0 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	18 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_Update/LOAD_next_pc1_135_Merge/merge_ack
      -- CP-element group 15: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_Update/LOAD_next_pc1_135_Merge/merge_req
      -- CP-element group 15: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_Update/LOAD_next_pc1_135_Merge/$exit
      -- CP-element group 15: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_Update/LOAD_next_pc1_135_Merge/$entry
      -- CP-element group 15: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_Update/word_access_complete/word_0/ca
      -- CP-element group 15: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_Update/word_access_complete/word_0/$exit
      -- CP-element group 15: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_Update/word_access_complete/$exit
      -- CP-element group 15: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_Update/$exit
      -- CP-element group 15: 	 assign_stmt_122_to_assign_stmt_136/LOAD_next_pc1_135_update_completed_
      -- 
    ca_676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_next_pc1_135_load_0_ack_1, ack => bz_CP_535_elements(15)); -- 
    -- CP-element group 16:  transition  delay-element  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	6 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	10 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_124_STORE_next_pc1_130_delay
      -- 
    -- Element group bz_CP_535_elements(16) is a control-delay.
    cp_element_16_delay: control_delay_element  generic map(name => " 16_delay", delay_value => 1)  port map(req => bz_CP_535_elements(6), ack => bz_CP_535_elements(16), clk => clk, reset =>reset);
    -- CP-element group 17:  transition  delay-element  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	13 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 assign_stmt_122_to_assign_stmt_136/STORE_next_pc1_130_LOAD_next_pc1_135_delay
      -- 
    -- Element group bz_CP_535_elements(17) is a control-delay.
    cp_element_17_delay: control_delay_element  generic map(name => " 17_delay", delay_value => 1)  port map(req => bz_CP_535_elements(11), ack => bz_CP_535_elements(17), clk => clk, reset =>reset);
    -- CP-element group 18:  join  transition  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	7 
    -- CP-element group 18: 	12 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 assign_stmt_122_to_assign_stmt_136/$exit
      -- CP-element group 18: 	 $exit
      -- 
    bz_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 22) := "bz_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= bz_CP_535_elements(7) & bz_CP_535_elements(12) & bz_CP_535_elements(15);
      gj_bz_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => bz_CP_535_elements(18), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u8_u8_127_wire : std_logic_vector(7 downto 0);
    signal LOAD_next_pc1_135_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_next_pc1_135_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_next_pc1_124_data_0 : std_logic_vector(7 downto 0);
    signal STORE_next_pc1_124_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_next_pc1_130_data_0 : std_logic_vector(7 downto 0);
    signal STORE_next_pc1_130_word_address_0 : std_logic_vector(0 downto 0);
    signal bzz_122 : std_logic_vector(31 downto 0);
    signal konst_126_wire_constant : std_logic_vector(7 downto 0);
    signal slice_132_wire : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    LOAD_next_pc1_135_word_address_0 <= "0";
    STORE_next_pc1_124_word_address_0 <= "0";
    STORE_next_pc1_130_word_address_0 <= "0";
    konst_126_wire_constant <= "00000001";
    slice_132_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      signal sample_req_ug, sample_ack_ug, update_req_ug, update_ack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      sample_req_ug(0) <= slice_132_inst_req_0;
      slice_132_inst_ack_0<= sample_ack_ug(0);
      update_req_ug(0) <= slice_132_inst_req_1;
      slice_132_inst_ack_1<= update_ack_ug(0);
      guard_vector(0) <=  not bzz_122(0);
      slice_132_inst_gI: SplitGuardInterface generic map(name => "slice_132_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_ug,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_ug,
        cr_in => update_req_ug,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_ug,
        guards => guard_vector); -- 
      slice_132_inst: SliceSplitProtocol generic map(name => "slice_132_inst", in_data_width => 32, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => rs2_data_buffer, dout => slice_132_wire, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_bzz_120_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_bzz_120_inst_req_0;
      W_bzz_120_inst_ack_0<= wack(0);
      rreq(0) <= W_bzz_120_inst_req_1;
      W_bzz_120_inst_ack_1<= rack(0);
      W_bzz_120_inst : InterlockBuffer generic map ( -- 
        name => "W_bzz_120_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rs1_data_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => bzz_122,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_next_pc1_135_gather_scatter
    process(LOAD_next_pc1_135_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_next_pc1_135_data_0;
      ov(7 downto 0) := iv;
      next_pc_buffer <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_next_pc1_124_gather_scatter
    process(ADD_u8_u8_127_wire) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u8_u8_127_wire;
      ov(7 downto 0) := iv;
      STORE_next_pc1_124_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_next_pc1_130_gather_scatter
    process(slice_132_wire) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := slice_132_wire;
      ov(7 downto 0) := iv;
      STORE_next_pc1_130_data_0 <= ov(7 downto 0);
      --
    end process;
    -- shared split operator group (0) : ADD_u8_u8_127_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pc_buffer;
      ADD_u8_u8_127_wire <= data_out(7 downto 0);
      guard_vector(0)  <= bzz_122(0);
      reqL_unguarded(0) <= ADD_u8_u8_127_inst_req_0;
      ADD_u8_u8_127_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_127_inst_req_1;
      ADD_u8_u8_127_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared load operator group (0) : LOAD_next_pc1_135_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_next_pc1_135_load_0_req_0;
      LOAD_next_pc1_135_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_next_pc1_135_load_0_req_1;
      LOAD_next_pc1_135_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_next_pc1_135_word_address_0;
      LOAD_next_pc1_135_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(0 downto 0),
          mtag => memory_space_1_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(7 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : STORE_next_pc1_130_store_0 STORE_next_pc1_124_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(1 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= STORE_next_pc1_130_store_0_req_0;
      reqL_unguarded(0) <= STORE_next_pc1_124_store_0_req_0;
      STORE_next_pc1_130_store_0_ack_0 <= ackL_unguarded(1);
      STORE_next_pc1_124_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= STORE_next_pc1_130_store_0_req_1;
      reqR_unguarded(0) <= STORE_next_pc1_124_store_0_req_1;
      STORE_next_pc1_130_store_0_ack_1 <= ackR_unguarded(1);
      STORE_next_pc1_124_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= bzz_122(0);
      guard_vector(1)  <=  not bzz_122(0);
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_next_pc1_130_word_address_0 & STORE_next_pc1_124_word_address_0;
      data_in <= STORE_next_pc1_130_data_0 & STORE_next_pc1_124_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(0 downto 0),
          mdata => memory_space_1_sr_data(7 downto 0),
          mtag => memory_space_1_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end bz_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity call is -- 
  generic (tag_length : integer); 
  port ( -- 
    rs1_data : in  std_logic_vector(31 downto 0);
    rs2_data : in  std_logic_vector(31 downto 0);
    rd : in  std_logic_vector(7 downto 0);
    pc : in  std_logic_vector(7 downto 0);
    next_pc : out  std_logic_vector(7 downto 0);
    accessreg_call_reqs : out  std_logic_vector(0 downto 0);
    accessreg_call_acks : in   std_logic_vector(0 downto 0);
    accessreg_call_data : out  std_logic_vector(40 downto 0);
    accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
    accessreg_return_reqs : out  std_logic_vector(0 downto 0);
    accessreg_return_acks : in   std_logic_vector(0 downto 0);
    accessreg_return_data : in   std_logic_vector(31 downto 0);
    accessreg_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity call;
architecture call_arch of call is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 80)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rs1_data_buffer :  std_logic_vector(31 downto 0);
  signal rs1_data_update_enable: Boolean;
  signal rs2_data_buffer :  std_logic_vector(31 downto 0);
  signal rs2_data_update_enable: Boolean;
  signal rd_buffer :  std_logic_vector(7 downto 0);
  signal rd_update_enable: Boolean;
  signal pc_buffer :  std_logic_vector(7 downto 0);
  signal pc_update_enable: Boolean;
  -- output port buffer signals
  signal next_pc_buffer :  std_logic_vector(7 downto 0);
  signal next_pc_update_enable: Boolean;
  signal call_CP_684_start: Boolean;
  signal call_CP_684_symbol: Boolean;
  -- volatile/operator module components. 
  component accessreg is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(7 downto 0);
      write_data : in  std_logic_vector(31 downto 0);
      read_data : out  std_logic_vector(31 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal CONCAT_u24_u32_151_inst_ack_1 : boolean;
  signal CONCAT_u24_u32_151_inst_req_1 : boolean;
  signal call_stmt_157_call_ack_1 : boolean;
  signal call_stmt_157_call_req_0 : boolean;
  signal call_stmt_157_call_req_1 : boolean;
  signal call_stmt_157_call_ack_0 : boolean;
  signal slice_160_inst_ack_1 : boolean;
  signal slice_160_inst_req_1 : boolean;
  signal slice_160_inst_ack_0 : boolean;
  signal CONCAT_u24_u32_151_inst_ack_0 : boolean;
  signal CONCAT_u24_u32_151_inst_req_0 : boolean;
  signal slice_160_inst_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "call_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 80) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= rs1_data;
  rs1_data_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= rs2_data;
  rs2_data_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(71 downto 64) <= rd;
  rd_buffer <= in_buffer_data_out(71 downto 64);
  in_buffer_data_in(79 downto 72) <= pc;
  pc_buffer <= in_buffer_data_out(79 downto 72);
  in_buffer_data_in(tag_length + 79 downto 80) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 79 downto 80);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  call_CP_684_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "call_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= next_pc_buffer;
  next_pc <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= call_CP_684_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= call_CP_684_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= call_CP_684_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  call_CP_684: Block -- control-path 
    signal call_CP_684_elements: BooleanArray(7 downto 0);
    -- 
  begin -- 
    call_CP_684_elements(0) <= call_CP_684_start;
    call_CP_684_symbol <= call_CP_684_elements(7);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0:  members (17) 
      -- CP-element group 0: 	 assign_stmt_152_to_assign_stmt_161/slice_160_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_152_to_assign_stmt_161/slice_160_update_start_
      -- CP-element group 0: 	 assign_stmt_152_to_assign_stmt_161/slice_160_sample_start_
      -- CP-element group 0: 	 assign_stmt_152_to_assign_stmt_161/CONCAT_u24_u32_151_Update/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_152_to_assign_stmt_161/slice_160_Update/$entry
      -- CP-element group 0: 	 assign_stmt_152_to_assign_stmt_161/call_stmt_157_Update/ccr
      -- CP-element group 0: 	 assign_stmt_152_to_assign_stmt_161/call_stmt_157_Update/$entry
      -- CP-element group 0: 	 assign_stmt_152_to_assign_stmt_161/CONCAT_u24_u32_151_Update/$entry
      -- CP-element group 0: 	 assign_stmt_152_to_assign_stmt_161/slice_160_Update/cr
      -- CP-element group 0: 	 assign_stmt_152_to_assign_stmt_161/call_stmt_157_update_start_
      -- CP-element group 0: 	 assign_stmt_152_to_assign_stmt_161/CONCAT_u24_u32_151_Sample/rr
      -- CP-element group 0: 	 assign_stmt_152_to_assign_stmt_161/CONCAT_u24_u32_151_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_152_to_assign_stmt_161/slice_160_Sample/rr
      -- CP-element group 0: 	 assign_stmt_152_to_assign_stmt_161/CONCAT_u24_u32_151_update_start_
      -- CP-element group 0: 	 assign_stmt_152_to_assign_stmt_161/CONCAT_u24_u32_151_sample_start_
      -- CP-element group 0: 	 assign_stmt_152_to_assign_stmt_161/$entry
      -- 
    rr_697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_CP_684_elements(0), ack => CONCAT_u24_u32_151_inst_req_0); -- 
    cr_702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_CP_684_elements(0), ack => CONCAT_u24_u32_151_inst_req_1); -- 
    ccr_716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_CP_684_elements(0), ack => call_stmt_157_call_req_1); -- 
    rr_725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_CP_684_elements(0), ack => slice_160_inst_req_0); -- 
    cr_730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_CP_684_elements(0), ack => slice_160_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_161/CONCAT_u24_u32_151_Sample/ra
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_161/CONCAT_u24_u32_151_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_152_to_assign_stmt_161/CONCAT_u24_u32_151_sample_completed_
      -- 
    ra_698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u24_u32_151_inst_ack_0, ack => call_CP_684_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_152_to_assign_stmt_161/CONCAT_u24_u32_151_Update/ca
      -- CP-element group 2: 	 assign_stmt_152_to_assign_stmt_161/call_stmt_157_Sample/crr
      -- CP-element group 2: 	 assign_stmt_152_to_assign_stmt_161/CONCAT_u24_u32_151_Update/$exit
      -- CP-element group 2: 	 assign_stmt_152_to_assign_stmt_161/call_stmt_157_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_152_to_assign_stmt_161/call_stmt_157_sample_start_
      -- CP-element group 2: 	 assign_stmt_152_to_assign_stmt_161/CONCAT_u24_u32_151_update_completed_
      -- 
    ca_703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u24_u32_151_inst_ack_1, ack => call_CP_684_elements(2)); -- 
    crr_711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_CP_684_elements(2), ack => call_stmt_157_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_152_to_assign_stmt_161/call_stmt_157_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_152_to_assign_stmt_161/call_stmt_157_Sample/cra
      -- CP-element group 3: 	 assign_stmt_152_to_assign_stmt_161/call_stmt_157_sample_completed_
      -- 
    cra_712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_157_call_ack_0, ack => call_CP_684_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_152_to_assign_stmt_161/call_stmt_157_Update/cca
      -- CP-element group 4: 	 assign_stmt_152_to_assign_stmt_161/call_stmt_157_Update/$exit
      -- CP-element group 4: 	 assign_stmt_152_to_assign_stmt_161/call_stmt_157_update_completed_
      -- 
    cca_717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_157_call_ack_1, ack => call_CP_684_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_152_to_assign_stmt_161/slice_160_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_152_to_assign_stmt_161/slice_160_sample_completed_
      -- CP-element group 5: 	 assign_stmt_152_to_assign_stmt_161/slice_160_Sample/ra
      -- 
    ra_726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_160_inst_ack_0, ack => call_CP_684_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_152_to_assign_stmt_161/slice_160_update_completed_
      -- CP-element group 6: 	 assign_stmt_152_to_assign_stmt_161/slice_160_Update/ca
      -- CP-element group 6: 	 assign_stmt_152_to_assign_stmt_161/slice_160_Update/$exit
      -- 
    ca_731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_160_inst_ack_1, ack => call_CP_684_elements(6)); -- 
    -- CP-element group 7:  join  transition  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 $exit
      -- CP-element group 7: 	 assign_stmt_152_to_assign_stmt_161/$exit
      -- 
    call_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 23) := "call_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= call_CP_684_elements(4) & call_CP_684_elements(6);
      gj_call_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => call_CP_684_elements(7), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_zero24_149_wire_constant : std_logic_vector(23 downto 0);
    signal dummy_157 : std_logic_vector(31 downto 0);
    signal konst_153_wire_constant : std_logic_vector(0 downto 0);
    signal pc_32_152 : std_logic_vector(31 downto 0);
    signal xxcallxxzero24 : std_logic_vector(23 downto 0);
    -- 
  begin -- 
    R_zero24_149_wire_constant <= "000000000000000000000000";
    konst_153_wire_constant <= "0";
    xxcallxxzero24 <= "000000000000000000000000";
    slice_160_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_160_inst_req_0;
      slice_160_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_160_inst_req_1;
      slice_160_inst_ack_1<= update_ack(0);
      slice_160_inst: SliceSplitProtocol generic map(name => "slice_160_inst", in_data_width => 32, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => rs1_data_buffer, dout => next_pc_buffer, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- shared split operator group (0) : CONCAT_u24_u32_151_inst 
    ApConcat_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_zero24_149_wire_constant & pc_buffer;
      pc_32_152 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u24_u32_151_inst_req_0;
      CONCAT_u24_u32_151_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u24_u32_151_inst_req_1;
      CONCAT_u24_u32_151_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_0_gI: SplitGuardInterface generic map(name => "ApConcat_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 24,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared call operator group (0) : call_stmt_157_call 
    accessreg_call_group_0: Block -- 
      signal data_in: std_logic_vector(40 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_157_call_req_0;
      call_stmt_157_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_157_call_req_1;
      call_stmt_157_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessreg_call_group_0_gI: SplitGuardInterface generic map(name => "accessreg_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_153_wire_constant & rd_buffer & pc_32_152;
      dummy_157 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 41,
        owidth => 41,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessreg_call_reqs(0),
          ackR => accessreg_call_acks(0),
          dataR => accessreg_call_data(40 downto 0),
          tagR => accessreg_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessreg_return_acks(0), -- cross-over
          ackL => accessreg_return_reqs(0), -- cross-over
          dataL => accessreg_return_data(31 downto 0),
          tagL => accessreg_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end call_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity cmp is -- 
  generic (tag_length : integer); 
  port ( -- 
    rs1_data : in  std_logic_vector(31 downto 0);
    rs2_data : in  std_logic_vector(31 downto 0);
    rd : in  std_logic_vector(7 downto 0);
    pc : in  std_logic_vector(7 downto 0);
    next_pc : out  std_logic_vector(7 downto 0);
    accessreg_call_reqs : out  std_logic_vector(0 downto 0);
    accessreg_call_acks : in   std_logic_vector(0 downto 0);
    accessreg_call_data : out  std_logic_vector(40 downto 0);
    accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
    accessreg_return_reqs : out  std_logic_vector(0 downto 0);
    accessreg_return_acks : in   std_logic_vector(0 downto 0);
    accessreg_return_data : in   std_logic_vector(31 downto 0);
    accessreg_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity cmp;
architecture cmp_arch of cmp is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 80)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rs1_data_buffer :  std_logic_vector(31 downto 0);
  signal rs1_data_update_enable: Boolean;
  signal rs2_data_buffer :  std_logic_vector(31 downto 0);
  signal rs2_data_update_enable: Boolean;
  signal rd_buffer :  std_logic_vector(7 downto 0);
  signal rd_update_enable: Boolean;
  signal pc_buffer :  std_logic_vector(7 downto 0);
  signal pc_update_enable: Boolean;
  -- output port buffer signals
  signal next_pc_buffer :  std_logic_vector(7 downto 0);
  signal next_pc_update_enable: Boolean;
  signal cmp_CP_732_start: Boolean;
  signal cmp_CP_732_symbol: Boolean;
  -- volatile/operator module components. 
  component accessreg is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(7 downto 0);
      write_data : in  std_logic_vector(31 downto 0);
      read_data : out  std_logic_vector(31 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal OR_u32_u32_189_inst_ack_1 : boolean;
  signal OR_u32_u32_189_inst_req_1 : boolean;
  signal ADD_u8_u8_199_inst_ack_0 : boolean;
  signal ADD_u8_u8_199_inst_req_0 : boolean;
  signal OR_u32_u32_189_inst_ack_0 : boolean;
  signal call_stmt_195_call_ack_1 : boolean;
  signal call_stmt_195_call_req_1 : boolean;
  signal call_stmt_195_call_ack_0 : boolean;
  signal call_stmt_195_call_req_0 : boolean;
  signal OR_u32_u32_189_inst_req_0 : boolean;
  signal ADD_u8_u8_199_inst_ack_1 : boolean;
  signal ADD_u8_u8_199_inst_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "cmp_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 80) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= rs1_data;
  rs1_data_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= rs2_data;
  rs2_data_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(71 downto 64) <= rd;
  rd_buffer <= in_buffer_data_out(71 downto 64);
  in_buffer_data_in(79 downto 72) <= pc;
  pc_buffer <= in_buffer_data_out(79 downto 72);
  in_buffer_data_in(tag_length + 79 downto 80) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 79 downto 80);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  cmp_CP_732_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "cmp_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= next_pc_buffer;
  next_pc <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= cmp_CP_732_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= cmp_CP_732_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= cmp_CP_732_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  cmp_CP_732: Block -- control-path 
    signal cmp_CP_732_elements: BooleanArray(7 downto 0);
    -- 
  begin -- 
    cmp_CP_732_elements(0) <= cmp_CP_732_start;
    cmp_CP_732_symbol <= cmp_CP_732_elements(7);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0:  members (17) 
      -- CP-element group 0: 	 assign_stmt_190_to_assign_stmt_200/$entry
      -- CP-element group 0: 	 assign_stmt_190_to_assign_stmt_200/OR_u32_u32_189_Update/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_190_to_assign_stmt_200/ADD_u8_u8_199_Sample/rr
      -- CP-element group 0: 	 assign_stmt_190_to_assign_stmt_200/ADD_u8_u8_199_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_190_to_assign_stmt_200/ADD_u8_u8_199_update_start_
      -- CP-element group 0: 	 assign_stmt_190_to_assign_stmt_200/ADD_u8_u8_199_sample_start_
      -- CP-element group 0: 	 assign_stmt_190_to_assign_stmt_200/OR_u32_u32_189_Update/$entry
      -- CP-element group 0: 	 assign_stmt_190_to_assign_stmt_200/call_stmt_195_update_start_
      -- CP-element group 0: 	 assign_stmt_190_to_assign_stmt_200/call_stmt_195_Update/ccr
      -- CP-element group 0: 	 assign_stmt_190_to_assign_stmt_200/call_stmt_195_Update/$entry
      -- CP-element group 0: 	 assign_stmt_190_to_assign_stmt_200/OR_u32_u32_189_Sample/rr
      -- CP-element group 0: 	 assign_stmt_190_to_assign_stmt_200/ADD_u8_u8_199_Update/cr
      -- CP-element group 0: 	 assign_stmt_190_to_assign_stmt_200/ADD_u8_u8_199_Update/$entry
      -- CP-element group 0: 	 assign_stmt_190_to_assign_stmt_200/OR_u32_u32_189_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_190_to_assign_stmt_200/OR_u32_u32_189_sample_start_
      -- CP-element group 0: 	 assign_stmt_190_to_assign_stmt_200/OR_u32_u32_189_update_start_
      -- 
    rr_745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => cmp_CP_732_elements(0), ack => OR_u32_u32_189_inst_req_0); -- 
    cr_750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => cmp_CP_732_elements(0), ack => OR_u32_u32_189_inst_req_1); -- 
    ccr_764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => cmp_CP_732_elements(0), ack => call_stmt_195_call_req_1); -- 
    rr_773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => cmp_CP_732_elements(0), ack => ADD_u8_u8_199_inst_req_0); -- 
    cr_778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => cmp_CP_732_elements(0), ack => ADD_u8_u8_199_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_190_to_assign_stmt_200/OR_u32_u32_189_Sample/ra
      -- CP-element group 1: 	 assign_stmt_190_to_assign_stmt_200/OR_u32_u32_189_sample_completed_
      -- CP-element group 1: 	 assign_stmt_190_to_assign_stmt_200/OR_u32_u32_189_Sample/$exit
      -- 
    ra_746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_189_inst_ack_0, ack => cmp_CP_732_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_190_to_assign_stmt_200/OR_u32_u32_189_update_completed_
      -- CP-element group 2: 	 assign_stmt_190_to_assign_stmt_200/OR_u32_u32_189_Update/ca
      -- CP-element group 2: 	 assign_stmt_190_to_assign_stmt_200/OR_u32_u32_189_Update/$exit
      -- CP-element group 2: 	 assign_stmt_190_to_assign_stmt_200/call_stmt_195_Sample/crr
      -- CP-element group 2: 	 assign_stmt_190_to_assign_stmt_200/call_stmt_195_sample_start_
      -- CP-element group 2: 	 assign_stmt_190_to_assign_stmt_200/call_stmt_195_Sample/$entry
      -- 
    ca_751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_189_inst_ack_1, ack => cmp_CP_732_elements(2)); -- 
    crr_759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => cmp_CP_732_elements(2), ack => call_stmt_195_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_190_to_assign_stmt_200/call_stmt_195_Sample/cra
      -- CP-element group 3: 	 assign_stmt_190_to_assign_stmt_200/call_stmt_195_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_190_to_assign_stmt_200/call_stmt_195_sample_completed_
      -- 
    cra_760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_195_call_ack_0, ack => cmp_CP_732_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_190_to_assign_stmt_200/call_stmt_195_update_completed_
      -- CP-element group 4: 	 assign_stmt_190_to_assign_stmt_200/call_stmt_195_Update/cca
      -- CP-element group 4: 	 assign_stmt_190_to_assign_stmt_200/call_stmt_195_Update/$exit
      -- 
    cca_765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_195_call_ack_1, ack => cmp_CP_732_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_190_to_assign_stmt_200/ADD_u8_u8_199_Sample/ra
      -- CP-element group 5: 	 assign_stmt_190_to_assign_stmt_200/ADD_u8_u8_199_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_190_to_assign_stmt_200/ADD_u8_u8_199_sample_completed_
      -- 
    ra_774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_199_inst_ack_0, ack => cmp_CP_732_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_190_to_assign_stmt_200/ADD_u8_u8_199_update_completed_
      -- CP-element group 6: 	 assign_stmt_190_to_assign_stmt_200/ADD_u8_u8_199_Update/ca
      -- CP-element group 6: 	 assign_stmt_190_to_assign_stmt_200/ADD_u8_u8_199_Update/$exit
      -- 
    ca_779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_199_inst_ack_1, ack => cmp_CP_732_elements(6)); -- 
    -- CP-element group 7:  join  transition  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 assign_stmt_190_to_assign_stmt_200/$exit
      -- CP-element group 7: 	 $exit
      -- 
    cmp_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 22) := "cmp_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= cmp_CP_732_elements(4) & cmp_CP_732_elements(6);
      gj_cmp_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => cmp_CP_732_elements(7), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u32_u1_172_wire : std_logic_vector(0 downto 0);
    signal MUX_175_wire : std_logic_vector(31 downto 0);
    signal MUX_181_wire : std_logic_vector(31 downto 0);
    signal MUX_188_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_182_wire : std_logic_vector(31 downto 0);
    signal UGT_u32_u1_185_wire : std_logic_vector(0 downto 0);
    signal ULT_u32_u1_178_wire : std_logic_vector(0 downto 0);
    signal dummy_195 : std_logic_vector(31 downto 0);
    signal konst_173_wire_constant : std_logic_vector(31 downto 0);
    signal konst_174_wire_constant : std_logic_vector(31 downto 0);
    signal konst_179_wire_constant : std_logic_vector(31 downto 0);
    signal konst_180_wire_constant : std_logic_vector(31 downto 0);
    signal konst_186_wire_constant : std_logic_vector(31 downto 0);
    signal konst_187_wire_constant : std_logic_vector(31 downto 0);
    signal konst_191_wire_constant : std_logic_vector(0 downto 0);
    signal konst_198_wire_constant : std_logic_vector(7 downto 0);
    signal output_190 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_173_wire_constant <= "00000000000000000000000000000000";
    konst_174_wire_constant <= "00000000000000000000000000000000";
    konst_179_wire_constant <= "11111111111111111111111111111111";
    konst_180_wire_constant <= "00000000000000000000000000000000";
    konst_186_wire_constant <= "00000000000000000000000000000001";
    konst_187_wire_constant <= "00000000000000000000000000000000";
    konst_191_wire_constant <= "0";
    konst_198_wire_constant <= "00000001";
    -- flow-through select operator MUX_175_inst
    MUX_175_wire <= konst_173_wire_constant when (EQ_u32_u1_172_wire(0) /=  '0') else konst_174_wire_constant;
    -- flow-through select operator MUX_181_inst
    MUX_181_wire <= konst_179_wire_constant when (ULT_u32_u1_178_wire(0) /=  '0') else konst_180_wire_constant;
    -- flow-through select operator MUX_188_inst
    MUX_188_wire <= konst_186_wire_constant when (UGT_u32_u1_185_wire(0) /=  '0') else konst_187_wire_constant;
    -- shared split operator group (0) : ADD_u8_u8_199_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pc_buffer;
      next_pc_buffer <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_199_inst_req_0;
      ADD_u8_u8_199_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_199_inst_req_1;
      ADD_u8_u8_199_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator EQ_u32_u1_172_inst
    process(rs1_data_buffer, rs2_data_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(rs1_data_buffer, rs2_data_buffer, tmp_var);
      EQ_u32_u1_172_wire <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_182_inst
    process(MUX_175_wire, MUX_181_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_175_wire, MUX_181_wire, tmp_var);
      OR_u32_u32_182_wire <= tmp_var; --
    end process;
    -- shared split operator group (3) : OR_u32_u32_189_inst 
    ApIntOr_group_3: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= OR_u32_u32_182_wire & MUX_188_wire;
      output_190 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_189_inst_req_0;
      OR_u32_u32_189_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_189_inst_req_1;
      OR_u32_u32_189_inst_ack_1 <= ackR_unguarded(0);
      ApIntOr_group_3_gI: SplitGuardInterface generic map(name => "ApIntOr_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- binary operator UGT_u32_u1_185_inst
    process(rs1_data_buffer, rs2_data_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(rs1_data_buffer, rs2_data_buffer, tmp_var);
      UGT_u32_u1_185_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_178_inst
    process(rs1_data_buffer, rs2_data_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(rs1_data_buffer, rs2_data_buffer, tmp_var);
      ULT_u32_u1_178_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_195_call 
    accessreg_call_group_0: Block -- 
      signal data_in: std_logic_vector(40 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_195_call_req_0;
      call_stmt_195_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_195_call_req_1;
      call_stmt_195_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessreg_call_group_0_gI: SplitGuardInterface generic map(name => "accessreg_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_191_wire_constant & rd_buffer & output_190;
      dummy_195 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 41,
        owidth => 41,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessreg_call_reqs(0),
          ackR => accessreg_call_acks(0),
          dataR => accessreg_call_data(40 downto 0),
          tagR => accessreg_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessreg_return_acks(0), -- cross-over
          ackL => accessreg_return_reqs(0), -- cross-over
          dataL => accessreg_return_data(31 downto 0),
          tagL => accessreg_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end cmp_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity halt is -- 
  generic (tag_length : integer); 
  port ( -- 
    pc : in  std_logic_vector(7 downto 0);
    next_pc : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity halt;
architecture halt_arch of halt is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal pc_buffer :  std_logic_vector(7 downto 0);
  signal pc_update_enable: Boolean;
  -- output port buffer signals
  signal next_pc_buffer :  std_logic_vector(7 downto 0);
  signal next_pc_update_enable: Boolean;
  signal halt_CP_783_start: Boolean;
  signal halt_CP_783_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ADD_u8_u8_211_inst_req_0 : boolean;
  signal ADD_u8_u8_211_inst_ack_0 : boolean;
  signal ADD_u8_u8_211_inst_req_1 : boolean;
  signal ADD_u8_u8_211_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "halt_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 8) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= pc;
  pc_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(tag_length + 7 downto 8) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 7 downto 8);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  halt_CP_783_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "halt_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= next_pc_buffer;
  next_pc <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= halt_CP_783_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= halt_CP_783_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= halt_CP_783_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  halt_CP_783: Block -- control-path 
    signal halt_CP_783_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    halt_CP_783_elements(0) <= halt_CP_783_start;
    halt_CP_783_symbol <= halt_CP_783_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_212/ADD_u8_u8_211_Sample/rr
      -- CP-element group 0: 	 assign_stmt_212/ADD_u8_u8_211_Update/$entry
      -- CP-element group 0: 	 assign_stmt_212/ADD_u8_u8_211_Update/cr
      -- CP-element group 0: 	 assign_stmt_212/$entry
      -- CP-element group 0: 	 assign_stmt_212/ADD_u8_u8_211_sample_start_
      -- CP-element group 0: 	 assign_stmt_212/ADD_u8_u8_211_update_start_
      -- CP-element group 0: 	 assign_stmt_212/ADD_u8_u8_211_Sample/$entry
      -- CP-element group 0: 	 $entry
      -- 
    rr_796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => halt_CP_783_elements(0), ack => ADD_u8_u8_211_inst_req_0); -- 
    cr_801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => halt_CP_783_elements(0), ack => ADD_u8_u8_211_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_212/ADD_u8_u8_211_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_212/ADD_u8_u8_211_Sample/ra
      -- CP-element group 1: 	 assign_stmt_212/ADD_u8_u8_211_sample_completed_
      -- 
    ra_797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_211_inst_ack_0, ack => halt_CP_783_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 assign_stmt_212/ADD_u8_u8_211_Update/$exit
      -- CP-element group 2: 	 assign_stmt_212/ADD_u8_u8_211_Update/ca
      -- CP-element group 2: 	 assign_stmt_212/$exit
      -- CP-element group 2: 	 assign_stmt_212/ADD_u8_u8_211_update_completed_
      -- CP-element group 2: 	 $exit
      -- 
    ca_802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_211_inst_ack_1, ack => halt_CP_783_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal konst_210_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_210_wire_constant <= "00000001";
    -- shared split operator group (0) : ADD_u8_u8_211_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pc_buffer;
      next_pc_buffer <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_211_inst_req_0;
      ADD_u8_u8_211_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_211_inst_req_1;
      ADD_u8_u8_211_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- 
  end Block; -- data_path
  -- 
end halt_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity init_mem is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(7 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity init_mem;
architecture init_mem_arch of init_mem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal init_mem_CP_803_start: Boolean;
  signal init_mem_CP_803_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_225_inst_req_0 : boolean;
  signal type_cast_225_inst_ack_0 : boolean;
  signal type_cast_225_inst_req_1 : boolean;
  signal type_cast_225_inst_ack_1 : boolean;
  signal array_obj_ref_228_store_0_req_0 : boolean;
  signal array_obj_ref_228_store_0_ack_0 : boolean;
  signal array_obj_ref_228_store_0_req_1 : boolean;
  signal array_obj_ref_228_store_0_ack_1 : boolean;
  signal ADD_u8_u8_234_inst_req_0 : boolean;
  signal ADD_u8_u8_234_inst_ack_0 : boolean;
  signal ADD_u8_u8_234_inst_req_1 : boolean;
  signal ADD_u8_u8_234_inst_ack_1 : boolean;
  signal if_stmt_236_branch_req_0 : boolean;
  signal if_stmt_236_branch_ack_1 : boolean;
  signal if_stmt_236_branch_ack_0 : boolean;
  signal phi_stmt_217_req_0 : boolean;
  signal NI_235_221_buf_req_0 : boolean;
  signal NI_235_221_buf_ack_0 : boolean;
  signal NI_235_221_buf_req_1 : boolean;
  signal NI_235_221_buf_ack_1 : boolean;
  signal phi_stmt_217_req_1 : boolean;
  signal phi_stmt_217_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "init_mem_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  init_mem_CP_803_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "init_mem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= init_mem_CP_803_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= init_mem_CP_803_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= init_mem_CP_803_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  init_mem_CP_803: Block -- control-path 
    signal init_mem_CP_803_elements: BooleanArray(16 downto 0);
    -- 
  begin -- 
    init_mem_CP_803_elements(0) <= init_mem_CP_803_start;
    init_mem_CP_803_symbol <= init_mem_CP_803_elements(10);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	11 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_215/$entry
      -- CP-element group 0: 	 branch_block_stmt_215/branch_block_stmt_215__entry__
      -- CP-element group 0: 	 branch_block_stmt_215/merge_stmt_216__entry__
      -- CP-element group 0: 	 branch_block_stmt_215/merge_stmt_216_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_215/merge_stmt_216__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_215/merge_stmt_216__entry___PhiReq/phi_stmt_217/$entry
      -- CP-element group 0: 	 branch_block_stmt_215/merge_stmt_216__entry___PhiReq/phi_stmt_217/phi_stmt_217_sources/$entry
      -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	16 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/type_cast_225_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/type_cast_225_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/type_cast_225_sample_completed_
      -- 
    ra_828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_225_inst_ack_0, ack => init_mem_CP_803_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	16 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/type_cast_225_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/type_cast_225_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/type_cast_225_update_completed_
      -- 
    ca_833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_225_inst_ack_1, ack => init_mem_CP_803_elements(2)); -- 
    -- CP-element group 3:  join  transition  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: 	16 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_Sample/array_obj_ref_228_Split/$entry
      -- CP-element group 3: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_Sample/array_obj_ref_228_Split/$exit
      -- CP-element group 3: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_Sample/array_obj_ref_228_Split/split_req
      -- CP-element group 3: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_Sample/array_obj_ref_228_Split/split_ack
      -- CP-element group 3: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_Sample/word_access_start/word_0/rr
      -- 
    rr_883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => init_mem_CP_803_elements(3), ack => array_obj_ref_228_store_0_req_0); -- 
    init_mem_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "init_mem_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= init_mem_CP_803_elements(2) & init_mem_CP_803_elements(16);
      gj_init_mem_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => init_mem_CP_803_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_Sample/word_access_start/$exit
      -- CP-element group 4: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_Sample/word_access_start/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_Sample/word_access_start/word_0/ra
      -- 
    ra_884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_228_store_0_ack_0, ack => init_mem_CP_803_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	16 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	8 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_Update/word_access_complete/$exit
      -- CP-element group 5: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_Update/word_access_complete/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_Update/word_access_complete/word_0/ca
      -- 
    ca_895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_228_store_0_ack_1, ack => init_mem_CP_803_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	16 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/ADD_u8_u8_234_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/ADD_u8_u8_234_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/ADD_u8_u8_234_Sample/ra
      -- 
    ra_904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_234_inst_ack_0, ack => init_mem_CP_803_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	16 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/ADD_u8_u8_234_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/ADD_u8_u8_234_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/ADD_u8_u8_234_Update/ca
      -- 
    ca_909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_234_inst_ack_1, ack => init_mem_CP_803_elements(7)); -- 
    -- CP-element group 8:  branch  join  transition  place  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	5 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: 	10 
    -- CP-element group 8:  members (24) 
      -- CP-element group 8: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235__exit__
      -- CP-element group 8: 	 branch_block_stmt_215/if_stmt_236__entry__
      -- CP-element group 8: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/$exit
      -- CP-element group 8: 	 branch_block_stmt_215/if_stmt_236_dead_link/$entry
      -- CP-element group 8: 	 branch_block_stmt_215/if_stmt_236_eval_test/$entry
      -- CP-element group 8: 	 branch_block_stmt_215/if_stmt_236_eval_test/$exit
      -- CP-element group 8: 	 branch_block_stmt_215/if_stmt_236_eval_test/ULT_u8_u1_239/$entry
      -- CP-element group 8: 	 branch_block_stmt_215/if_stmt_236_eval_test/ULT_u8_u1_239/$exit
      -- CP-element group 8: 	 branch_block_stmt_215/if_stmt_236_eval_test/ULT_u8_u1_239/ULT_u8_u1_239_inputs/$entry
      -- CP-element group 8: 	 branch_block_stmt_215/if_stmt_236_eval_test/ULT_u8_u1_239/ULT_u8_u1_239_inputs/$exit
      -- CP-element group 8: 	 branch_block_stmt_215/if_stmt_236_eval_test/ULT_u8_u1_239/SplitProtocol/$entry
      -- CP-element group 8: 	 branch_block_stmt_215/if_stmt_236_eval_test/ULT_u8_u1_239/SplitProtocol/$exit
      -- CP-element group 8: 	 branch_block_stmt_215/if_stmt_236_eval_test/ULT_u8_u1_239/SplitProtocol/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_215/if_stmt_236_eval_test/ULT_u8_u1_239/SplitProtocol/Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_215/if_stmt_236_eval_test/ULT_u8_u1_239/SplitProtocol/Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_215/if_stmt_236_eval_test/ULT_u8_u1_239/SplitProtocol/Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_215/if_stmt_236_eval_test/ULT_u8_u1_239/SplitProtocol/Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_215/if_stmt_236_eval_test/ULT_u8_u1_239/SplitProtocol/Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_215/if_stmt_236_eval_test/ULT_u8_u1_239/SplitProtocol/Update/cr
      -- CP-element group 8: 	 branch_block_stmt_215/if_stmt_236_eval_test/ULT_u8_u1_239/SplitProtocol/Update/ca
      -- CP-element group 8: 	 branch_block_stmt_215/if_stmt_236_eval_test/branch_req
      -- CP-element group 8: 	 branch_block_stmt_215/ULT_u8_u1_239_place
      -- CP-element group 8: 	 branch_block_stmt_215/if_stmt_236_if_link/$entry
      -- CP-element group 8: 	 branch_block_stmt_215/if_stmt_236_else_link/$entry
      -- 
    branch_req_936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => init_mem_CP_803_elements(8), ack => if_stmt_236_branch_req_0); -- 
    init_mem_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "init_mem_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= init_mem_CP_803_elements(5) & init_mem_CP_803_elements(7);
      gj_init_mem_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => init_mem_CP_803_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  fork  transition  place  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9:  members (11) 
      -- CP-element group 9: 	 branch_block_stmt_215/if_stmt_236_if_link/$exit
      -- CP-element group 9: 	 branch_block_stmt_215/if_stmt_236_if_link/if_choice_transition
      -- CP-element group 9: 	 branch_block_stmt_215/loopback
      -- CP-element group 9: 	 branch_block_stmt_215/loopback_PhiReq/$entry
      -- CP-element group 9: 	 branch_block_stmt_215/loopback_PhiReq/phi_stmt_217/$entry
      -- CP-element group 9: 	 branch_block_stmt_215/loopback_PhiReq/phi_stmt_217/phi_stmt_217_sources/$entry
      -- CP-element group 9: 	 branch_block_stmt_215/loopback_PhiReq/phi_stmt_217/phi_stmt_217_sources/Interlock/$entry
      -- CP-element group 9: 	 branch_block_stmt_215/loopback_PhiReq/phi_stmt_217/phi_stmt_217_sources/Interlock/Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_215/loopback_PhiReq/phi_stmt_217/phi_stmt_217_sources/Interlock/Sample/req
      -- CP-element group 9: 	 branch_block_stmt_215/loopback_PhiReq/phi_stmt_217/phi_stmt_217_sources/Interlock/Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_215/loopback_PhiReq/phi_stmt_217/phi_stmt_217_sources/Interlock/Update/req
      -- 
    if_choice_transition_941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_236_branch_ack_1, ack => init_mem_CP_803_elements(9)); -- 
    req_977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => init_mem_CP_803_elements(9), ack => NI_235_221_buf_req_0); -- 
    req_982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => init_mem_CP_803_elements(9), ack => NI_235_221_buf_req_1); -- 
    -- CP-element group 10:  merge  transition  place  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 $exit
      -- CP-element group 10: 	 branch_block_stmt_215/$exit
      -- CP-element group 10: 	 branch_block_stmt_215/branch_block_stmt_215__exit__
      -- CP-element group 10: 	 branch_block_stmt_215/if_stmt_236__exit__
      -- CP-element group 10: 	 branch_block_stmt_215/if_stmt_236_else_link/$exit
      -- CP-element group 10: 	 branch_block_stmt_215/if_stmt_236_else_link/else_choice_transition
      -- 
    else_choice_transition_945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_236_branch_ack_0, ack => init_mem_CP_803_elements(10)); -- 
    -- CP-element group 11:  transition  output  delay-element  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	15 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_215/merge_stmt_216__entry___PhiReq/$exit
      -- CP-element group 11: 	 branch_block_stmt_215/merge_stmt_216__entry___PhiReq/phi_stmt_217/$exit
      -- CP-element group 11: 	 branch_block_stmt_215/merge_stmt_216__entry___PhiReq/phi_stmt_217/phi_stmt_217_sources/$exit
      -- CP-element group 11: 	 branch_block_stmt_215/merge_stmt_216__entry___PhiReq/phi_stmt_217/phi_stmt_217_sources/type_cast_220_konst_delay_trans
      -- CP-element group 11: 	 branch_block_stmt_215/merge_stmt_216__entry___PhiReq/phi_stmt_217/phi_stmt_217_req
      -- 
    phi_stmt_217_req_961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_217_req_961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => init_mem_CP_803_elements(11), ack => phi_stmt_217_req_0); -- 
    -- Element group init_mem_CP_803_elements(11) is a control-delay.
    cp_element_11_delay: control_delay_element  generic map(name => " 11_delay", delay_value => 1)  port map(req => init_mem_CP_803_elements(0), ack => init_mem_CP_803_elements(11), clk => clk, reset =>reset);
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_215/loopback_PhiReq/phi_stmt_217/phi_stmt_217_sources/Interlock/Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_215/loopback_PhiReq/phi_stmt_217/phi_stmt_217_sources/Interlock/Sample/ack
      -- 
    ack_978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NI_235_221_buf_ack_0, ack => init_mem_CP_803_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_215/loopback_PhiReq/phi_stmt_217/phi_stmt_217_sources/Interlock/Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_215/loopback_PhiReq/phi_stmt_217/phi_stmt_217_sources/Interlock/Update/ack
      -- 
    ack_983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NI_235_221_buf_ack_1, ack => init_mem_CP_803_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (5) 
      -- CP-element group 14: 	 branch_block_stmt_215/loopback_PhiReq/$exit
      -- CP-element group 14: 	 branch_block_stmt_215/loopback_PhiReq/phi_stmt_217/$exit
      -- CP-element group 14: 	 branch_block_stmt_215/loopback_PhiReq/phi_stmt_217/phi_stmt_217_sources/$exit
      -- CP-element group 14: 	 branch_block_stmt_215/loopback_PhiReq/phi_stmt_217/phi_stmt_217_sources/Interlock/$exit
      -- CP-element group 14: 	 branch_block_stmt_215/loopback_PhiReq/phi_stmt_217/phi_stmt_217_req
      -- 
    phi_stmt_217_req_984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_217_req_984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => init_mem_CP_803_elements(14), ack => phi_stmt_217_req_1); -- 
    init_mem_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "init_mem_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= init_mem_CP_803_elements(12) & init_mem_CP_803_elements(13);
      gj_init_mem_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => init_mem_CP_803_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  merge  transition  place  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	11 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_215/merge_stmt_216_PhiReqMerge
      -- CP-element group 15: 	 branch_block_stmt_215/merge_stmt_216_PhiAck/$entry
      -- 
    init_mem_CP_803_elements(15) <= OrReduce(init_mem_CP_803_elements(11) & init_mem_CP_803_elements(14));
    -- CP-element group 16:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	1 
    -- CP-element group 16: 	2 
    -- CP-element group 16: 	3 
    -- CP-element group 16: 	5 
    -- CP-element group 16: 	6 
    -- CP-element group 16: 	7 
    -- CP-element group 16:  members (48) 
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/type_cast_225_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/type_cast_225_Sample/rr
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/type_cast_225_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/type_cast_225_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_update_start_
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_word_address_calculated
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_root_address_calculated
      -- CP-element group 16: 	 branch_block_stmt_215/merge_stmt_216__exit__
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235__entry__
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/$entry
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/type_cast_225_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/type_cast_225_update_start_
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_offset_calculated
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_index_resized_0
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_index_scaled_0
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_index_computed_0
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_index_resize_0/$entry
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_index_resize_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_index_resize_0/index_resize_req
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_index_resize_0/index_resize_ack
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_index_scale_0/$entry
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_index_scale_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_index_scale_0/scale_rename_req
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_index_scale_0/scale_rename_ack
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_final_index_sum_regn/$entry
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_final_index_sum_regn/$exit
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_final_index_sum_regn/req
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_final_index_sum_regn/ack
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_base_plus_offset/$entry
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_base_plus_offset/$exit
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_base_plus_offset/sum_rename_req
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_base_plus_offset/sum_rename_ack
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_word_addrgen/$entry
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_word_addrgen/$exit
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_word_addrgen/root_register_req
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_word_addrgen/root_register_ack
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_Update/word_access_complete/$entry
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_Update/word_access_complete/word_0/$entry
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/array_obj_ref_228_Update/word_access_complete/word_0/cr
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/ADD_u8_u8_234_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/ADD_u8_u8_234_update_start_
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/ADD_u8_u8_234_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/ADD_u8_u8_234_Sample/rr
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/ADD_u8_u8_234_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_215/assign_stmt_226_to_assign_stmt_235/ADD_u8_u8_234_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_215/merge_stmt_216_PhiAck/$exit
      -- CP-element group 16: 	 branch_block_stmt_215/merge_stmt_216_PhiAck/phi_stmt_217_ack
      -- 
    phi_stmt_217_ack_989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_217_ack_0, ack => init_mem_CP_803_elements(16)); -- 
    rr_827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => init_mem_CP_803_elements(16), ack => type_cast_225_inst_req_0); -- 
    cr_832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => init_mem_CP_803_elements(16), ack => type_cast_225_inst_req_1); -- 
    cr_894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => init_mem_CP_803_elements(16), ack => array_obj_ref_228_store_0_req_1); -- 
    rr_903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => init_mem_CP_803_elements(16), ack => ADD_u8_u8_234_inst_req_0); -- 
    cr_908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => init_mem_CP_803_elements(16), ack => ADD_u8_u8_234_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal I_217 : std_logic_vector(7 downto 0);
    signal NII_226 : std_logic_vector(31 downto 0);
    signal NI_235 : std_logic_vector(7 downto 0);
    signal NI_235_221_buffered : std_logic_vector(7 downto 0);
    signal R_I_227_resized : std_logic_vector(7 downto 0);
    signal R_I_227_scaled : std_logic_vector(7 downto 0);
    signal ULT_u8_u1_239_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_228_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_228_final_offset : std_logic_vector(7 downto 0);
    signal array_obj_ref_228_offset_scale_factor_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_228_resized_base_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_228_root_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_228_word_address_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_228_word_offset_0 : std_logic_vector(7 downto 0);
    signal konst_233_wire_constant : std_logic_vector(7 downto 0);
    signal konst_238_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_220_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_228_offset_scale_factor_0 <= "00000001";
    array_obj_ref_228_resized_base_address <= "00000000";
    array_obj_ref_228_word_offset_0 <= "00000000";
    konst_233_wire_constant <= "00000001";
    konst_238_wire_constant <= "00001010";
    type_cast_220_wire_constant <= "00000000";
    phi_stmt_217: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_220_wire_constant & NI_235_221_buffered;
      req <= phi_stmt_217_req_0 & phi_stmt_217_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_217",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_217_ack_0,
          idata => idata,
          odata => I_217,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_217
    NI_235_221_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= NI_235_221_buf_req_0;
      NI_235_221_buf_ack_0<= wack(0);
      rreq(0) <= NI_235_221_buf_req_1;
      NI_235_221_buf_ack_1<= rack(0);
      NI_235_221_buf : InterlockBuffer generic map ( -- 
        name => "NI_235_221_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => NI_235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NI_235_221_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_225_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_225_inst_req_0;
      type_cast_225_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_225_inst_req_1;
      type_cast_225_inst_ack_1<= rack(0);
      type_cast_225_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_225_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => I_217,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NII_226,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_228_addr_0
    process(array_obj_ref_228_root_address) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_228_root_address;
      ov(7 downto 0) := iv;
      array_obj_ref_228_word_address_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_228_gather_scatter
    process(NII_226) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := NII_226;
      ov(31 downto 0) := iv;
      array_obj_ref_228_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_228_index_0_rename
    process(R_I_227_resized) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_I_227_resized;
      ov(7 downto 0) := iv;
      R_I_227_scaled <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_228_index_0_resize
    process(I_217) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_217;
      ov(7 downto 0) := iv;
      R_I_227_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_228_index_offset
    process(R_I_227_scaled) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_I_227_scaled;
      ov(7 downto 0) := iv;
      array_obj_ref_228_final_offset <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_228_root_address_inst
    process(array_obj_ref_228_final_offset) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_228_final_offset;
      ov(7 downto 0) := iv;
      array_obj_ref_228_root_address <= ov(7 downto 0);
      --
    end process;
    if_stmt_236_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u8_u1_239_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_236_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_236_branch_req_0,
          ack0 => if_stmt_236_branch_ack_0,
          ack1 => if_stmt_236_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u8_u8_234_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= I_217;
      NI_235 <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_234_inst_req_0;
      ADD_u8_u8_234_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_234_inst_req_1;
      ADD_u8_u8_234_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator ULT_u8_u1_239_inst
    process(I_217) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(I_217, konst_238_wire_constant, tmp_var);
      ULT_u8_u1_239_wire <= tmp_var; --
    end process;
    -- shared store operator group (0) : array_obj_ref_228_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(7 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_228_store_0_req_0;
      array_obj_ref_228_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_228_store_0_req_1;
      array_obj_ref_228_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_228_word_address_0;
      data_in <= array_obj_ref_228_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 8,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(7 downto 0),
          mdata => memory_space_0_sr_data(31 downto 0),
          mtag => memory_space_0_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end init_mem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity init_reg is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(7 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity init_reg;
architecture init_reg_arch of init_reg is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal init_reg_CP_990_start: Boolean;
  signal init_reg_CP_990_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_255_inst_req_0 : boolean;
  signal type_cast_255_inst_ack_0 : boolean;
  signal type_cast_255_inst_req_1 : boolean;
  signal type_cast_255_inst_ack_1 : boolean;
  signal array_obj_ref_258_store_0_req_0 : boolean;
  signal array_obj_ref_258_store_0_ack_0 : boolean;
  signal array_obj_ref_258_store_0_req_1 : boolean;
  signal array_obj_ref_258_store_0_ack_1 : boolean;
  signal ADD_u8_u8_264_inst_req_0 : boolean;
  signal ADD_u8_u8_264_inst_ack_0 : boolean;
  signal ADD_u8_u8_264_inst_req_1 : boolean;
  signal ADD_u8_u8_264_inst_ack_1 : boolean;
  signal if_stmt_266_branch_req_0 : boolean;
  signal if_stmt_266_branch_ack_1 : boolean;
  signal if_stmt_266_branch_ack_0 : boolean;
  signal phi_stmt_247_req_0 : boolean;
  signal NJ_265_251_buf_req_0 : boolean;
  signal NJ_265_251_buf_ack_0 : boolean;
  signal NJ_265_251_buf_req_1 : boolean;
  signal NJ_265_251_buf_ack_1 : boolean;
  signal phi_stmt_247_req_1 : boolean;
  signal phi_stmt_247_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "init_reg_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  init_reg_CP_990_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "init_reg_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= init_reg_CP_990_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= init_reg_CP_990_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= init_reg_CP_990_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  init_reg_CP_990: Block -- control-path 
    signal init_reg_CP_990_elements: BooleanArray(16 downto 0);
    -- 
  begin -- 
    init_reg_CP_990_elements(0) <= init_reg_CP_990_start;
    init_reg_CP_990_symbol <= init_reg_CP_990_elements(10);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	11 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_245/$entry
      -- CP-element group 0: 	 branch_block_stmt_245/branch_block_stmt_245__entry__
      -- CP-element group 0: 	 branch_block_stmt_245/merge_stmt_246__entry__
      -- CP-element group 0: 	 branch_block_stmt_245/merge_stmt_246_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_245/merge_stmt_246__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_245/merge_stmt_246__entry___PhiReq/phi_stmt_247/$entry
      -- CP-element group 0: 	 branch_block_stmt_245/merge_stmt_246__entry___PhiReq/phi_stmt_247/phi_stmt_247_sources/$entry
      -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	16 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/type_cast_255_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/type_cast_255_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/type_cast_255_Sample/ra
      -- 
    ra_1015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_255_inst_ack_0, ack => init_reg_CP_990_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	16 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/type_cast_255_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/type_cast_255_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/type_cast_255_Update/ca
      -- 
    ca_1020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_255_inst_ack_1, ack => init_reg_CP_990_elements(2)); -- 
    -- CP-element group 3:  join  transition  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: 	16 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_Sample/array_obj_ref_258_Split/$entry
      -- CP-element group 3: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_Sample/array_obj_ref_258_Split/$exit
      -- CP-element group 3: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_Sample/array_obj_ref_258_Split/split_req
      -- CP-element group 3: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_Sample/array_obj_ref_258_Split/split_ack
      -- CP-element group 3: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_Sample/word_access_start/$entry
      -- CP-element group 3: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_Sample/word_access_start/word_0/rr
      -- 
    rr_1070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => init_reg_CP_990_elements(3), ack => array_obj_ref_258_store_0_req_0); -- 
    init_reg_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "init_reg_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= init_reg_CP_990_elements(2) & init_reg_CP_990_elements(16);
      gj_init_reg_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => init_reg_CP_990_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_Sample/word_access_start/$exit
      -- CP-element group 4: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_Sample/word_access_start/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_Sample/word_access_start/word_0/ra
      -- 
    ra_1071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_258_store_0_ack_0, ack => init_reg_CP_990_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	16 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	8 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_Update/word_access_complete/$exit
      -- CP-element group 5: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_Update/word_access_complete/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_Update/word_access_complete/word_0/ca
      -- 
    ca_1082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_258_store_0_ack_1, ack => init_reg_CP_990_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	16 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/ADD_u8_u8_264_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/ADD_u8_u8_264_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/ADD_u8_u8_264_Sample/ra
      -- 
    ra_1091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_264_inst_ack_0, ack => init_reg_CP_990_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	16 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/ADD_u8_u8_264_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/ADD_u8_u8_264_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/ADD_u8_u8_264_Update/ca
      -- 
    ca_1096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_264_inst_ack_1, ack => init_reg_CP_990_elements(7)); -- 
    -- CP-element group 8:  branch  join  transition  place  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	5 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: 	10 
    -- CP-element group 8:  members (24) 
      -- CP-element group 8: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265__exit__
      -- CP-element group 8: 	 branch_block_stmt_245/if_stmt_266__entry__
      -- CP-element group 8: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/$exit
      -- CP-element group 8: 	 branch_block_stmt_245/if_stmt_266_dead_link/$entry
      -- CP-element group 8: 	 branch_block_stmt_245/if_stmt_266_eval_test/$entry
      -- CP-element group 8: 	 branch_block_stmt_245/if_stmt_266_eval_test/$exit
      -- CP-element group 8: 	 branch_block_stmt_245/if_stmt_266_eval_test/ULT_u8_u1_269/$entry
      -- CP-element group 8: 	 branch_block_stmt_245/if_stmt_266_eval_test/ULT_u8_u1_269/$exit
      -- CP-element group 8: 	 branch_block_stmt_245/if_stmt_266_eval_test/ULT_u8_u1_269/ULT_u8_u1_269_inputs/$entry
      -- CP-element group 8: 	 branch_block_stmt_245/if_stmt_266_eval_test/ULT_u8_u1_269/ULT_u8_u1_269_inputs/$exit
      -- CP-element group 8: 	 branch_block_stmt_245/if_stmt_266_eval_test/ULT_u8_u1_269/SplitProtocol/$entry
      -- CP-element group 8: 	 branch_block_stmt_245/if_stmt_266_eval_test/ULT_u8_u1_269/SplitProtocol/$exit
      -- CP-element group 8: 	 branch_block_stmt_245/if_stmt_266_eval_test/ULT_u8_u1_269/SplitProtocol/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_245/if_stmt_266_eval_test/ULT_u8_u1_269/SplitProtocol/Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_245/if_stmt_266_eval_test/ULT_u8_u1_269/SplitProtocol/Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_245/if_stmt_266_eval_test/ULT_u8_u1_269/SplitProtocol/Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_245/if_stmt_266_eval_test/ULT_u8_u1_269/SplitProtocol/Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_245/if_stmt_266_eval_test/ULT_u8_u1_269/SplitProtocol/Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_245/if_stmt_266_eval_test/ULT_u8_u1_269/SplitProtocol/Update/cr
      -- CP-element group 8: 	 branch_block_stmt_245/if_stmt_266_eval_test/ULT_u8_u1_269/SplitProtocol/Update/ca
      -- CP-element group 8: 	 branch_block_stmt_245/if_stmt_266_eval_test/branch_req
      -- CP-element group 8: 	 branch_block_stmt_245/ULT_u8_u1_269_place
      -- CP-element group 8: 	 branch_block_stmt_245/if_stmt_266_if_link/$entry
      -- CP-element group 8: 	 branch_block_stmt_245/if_stmt_266_else_link/$entry
      -- 
    branch_req_1123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => init_reg_CP_990_elements(8), ack => if_stmt_266_branch_req_0); -- 
    init_reg_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "init_reg_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= init_reg_CP_990_elements(5) & init_reg_CP_990_elements(7);
      gj_init_reg_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => init_reg_CP_990_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  fork  transition  place  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9:  members (11) 
      -- CP-element group 9: 	 branch_block_stmt_245/if_stmt_266_if_link/$exit
      -- CP-element group 9: 	 branch_block_stmt_245/if_stmt_266_if_link/if_choice_transition
      -- CP-element group 9: 	 branch_block_stmt_245/loopback
      -- CP-element group 9: 	 branch_block_stmt_245/loopback_PhiReq/$entry
      -- CP-element group 9: 	 branch_block_stmt_245/loopback_PhiReq/phi_stmt_247/$entry
      -- CP-element group 9: 	 branch_block_stmt_245/loopback_PhiReq/phi_stmt_247/phi_stmt_247_sources/$entry
      -- CP-element group 9: 	 branch_block_stmt_245/loopback_PhiReq/phi_stmt_247/phi_stmt_247_sources/Interlock/$entry
      -- CP-element group 9: 	 branch_block_stmt_245/loopback_PhiReq/phi_stmt_247/phi_stmt_247_sources/Interlock/Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_245/loopback_PhiReq/phi_stmt_247/phi_stmt_247_sources/Interlock/Sample/req
      -- CP-element group 9: 	 branch_block_stmt_245/loopback_PhiReq/phi_stmt_247/phi_stmt_247_sources/Interlock/Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_245/loopback_PhiReq/phi_stmt_247/phi_stmt_247_sources/Interlock/Update/req
      -- 
    if_choice_transition_1128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_266_branch_ack_1, ack => init_reg_CP_990_elements(9)); -- 
    req_1164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => init_reg_CP_990_elements(9), ack => NJ_265_251_buf_req_0); -- 
    req_1169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => init_reg_CP_990_elements(9), ack => NJ_265_251_buf_req_1); -- 
    -- CP-element group 10:  merge  transition  place  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 $exit
      -- CP-element group 10: 	 branch_block_stmt_245/$exit
      -- CP-element group 10: 	 branch_block_stmt_245/branch_block_stmt_245__exit__
      -- CP-element group 10: 	 branch_block_stmt_245/if_stmt_266__exit__
      -- CP-element group 10: 	 branch_block_stmt_245/if_stmt_266_else_link/$exit
      -- CP-element group 10: 	 branch_block_stmt_245/if_stmt_266_else_link/else_choice_transition
      -- 
    else_choice_transition_1132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_266_branch_ack_0, ack => init_reg_CP_990_elements(10)); -- 
    -- CP-element group 11:  transition  output  delay-element  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	15 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_245/merge_stmt_246__entry___PhiReq/$exit
      -- CP-element group 11: 	 branch_block_stmt_245/merge_stmt_246__entry___PhiReq/phi_stmt_247/$exit
      -- CP-element group 11: 	 branch_block_stmt_245/merge_stmt_246__entry___PhiReq/phi_stmt_247/phi_stmt_247_sources/$exit
      -- CP-element group 11: 	 branch_block_stmt_245/merge_stmt_246__entry___PhiReq/phi_stmt_247/phi_stmt_247_sources/type_cast_250_konst_delay_trans
      -- CP-element group 11: 	 branch_block_stmt_245/merge_stmt_246__entry___PhiReq/phi_stmt_247/phi_stmt_247_req
      -- 
    phi_stmt_247_req_1148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_247_req_1148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => init_reg_CP_990_elements(11), ack => phi_stmt_247_req_0); -- 
    -- Element group init_reg_CP_990_elements(11) is a control-delay.
    cp_element_11_delay: control_delay_element  generic map(name => " 11_delay", delay_value => 1)  port map(req => init_reg_CP_990_elements(0), ack => init_reg_CP_990_elements(11), clk => clk, reset =>reset);
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_245/loopback_PhiReq/phi_stmt_247/phi_stmt_247_sources/Interlock/Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_245/loopback_PhiReq/phi_stmt_247/phi_stmt_247_sources/Interlock/Sample/ack
      -- 
    ack_1165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NJ_265_251_buf_ack_0, ack => init_reg_CP_990_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_245/loopback_PhiReq/phi_stmt_247/phi_stmt_247_sources/Interlock/Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_245/loopback_PhiReq/phi_stmt_247/phi_stmt_247_sources/Interlock/Update/ack
      -- 
    ack_1170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NJ_265_251_buf_ack_1, ack => init_reg_CP_990_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (5) 
      -- CP-element group 14: 	 branch_block_stmt_245/loopback_PhiReq/$exit
      -- CP-element group 14: 	 branch_block_stmt_245/loopback_PhiReq/phi_stmt_247/$exit
      -- CP-element group 14: 	 branch_block_stmt_245/loopback_PhiReq/phi_stmt_247/phi_stmt_247_sources/$exit
      -- CP-element group 14: 	 branch_block_stmt_245/loopback_PhiReq/phi_stmt_247/phi_stmt_247_sources/Interlock/$exit
      -- CP-element group 14: 	 branch_block_stmt_245/loopback_PhiReq/phi_stmt_247/phi_stmt_247_req
      -- 
    phi_stmt_247_req_1171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_247_req_1171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => init_reg_CP_990_elements(14), ack => phi_stmt_247_req_1); -- 
    init_reg_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "init_reg_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= init_reg_CP_990_elements(12) & init_reg_CP_990_elements(13);
      gj_init_reg_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => init_reg_CP_990_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  merge  transition  place  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	11 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_245/merge_stmt_246_PhiReqMerge
      -- CP-element group 15: 	 branch_block_stmt_245/merge_stmt_246_PhiAck/$entry
      -- 
    init_reg_CP_990_elements(15) <= OrReduce(init_reg_CP_990_elements(11) & init_reg_CP_990_elements(14));
    -- CP-element group 16:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	1 
    -- CP-element group 16: 	2 
    -- CP-element group 16: 	3 
    -- CP-element group 16: 	5 
    -- CP-element group 16: 	6 
    -- CP-element group 16: 	7 
    -- CP-element group 16:  members (48) 
      -- CP-element group 16: 	 branch_block_stmt_245/merge_stmt_246__exit__
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265__entry__
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/$entry
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/type_cast_255_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/type_cast_255_update_start_
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/type_cast_255_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/type_cast_255_Sample/rr
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/type_cast_255_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/type_cast_255_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_update_start_
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_word_address_calculated
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_root_address_calculated
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_offset_calculated
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_index_resized_0
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_index_scaled_0
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_index_computed_0
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_index_resize_0/$entry
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_index_resize_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_index_resize_0/index_resize_req
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_index_resize_0/index_resize_ack
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_index_scale_0/$entry
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_index_scale_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_index_scale_0/scale_rename_req
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_index_scale_0/scale_rename_ack
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_final_index_sum_regn/$entry
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_final_index_sum_regn/$exit
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_final_index_sum_regn/req
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_final_index_sum_regn/ack
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_base_plus_offset/$entry
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_base_plus_offset/$exit
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_base_plus_offset/sum_rename_req
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_base_plus_offset/sum_rename_ack
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_word_addrgen/$entry
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_word_addrgen/$exit
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_word_addrgen/root_register_req
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_word_addrgen/root_register_ack
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_Update/word_access_complete/$entry
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_Update/word_access_complete/word_0/$entry
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/array_obj_ref_258_Update/word_access_complete/word_0/cr
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/ADD_u8_u8_264_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/ADD_u8_u8_264_update_start_
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/ADD_u8_u8_264_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/ADD_u8_u8_264_Sample/rr
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/ADD_u8_u8_264_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_245/assign_stmt_256_to_assign_stmt_265/ADD_u8_u8_264_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_245/merge_stmt_246_PhiAck/$exit
      -- CP-element group 16: 	 branch_block_stmt_245/merge_stmt_246_PhiAck/phi_stmt_247_ack
      -- 
    phi_stmt_247_ack_1176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_247_ack_0, ack => init_reg_CP_990_elements(16)); -- 
    rr_1014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => init_reg_CP_990_elements(16), ack => type_cast_255_inst_req_0); -- 
    cr_1019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => init_reg_CP_990_elements(16), ack => type_cast_255_inst_req_1); -- 
    cr_1081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => init_reg_CP_990_elements(16), ack => array_obj_ref_258_store_0_req_1); -- 
    rr_1090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => init_reg_CP_990_elements(16), ack => ADD_u8_u8_264_inst_req_0); -- 
    cr_1095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => init_reg_CP_990_elements(16), ack => ADD_u8_u8_264_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal J_247 : std_logic_vector(7 downto 0);
    signal NJJ_256 : std_logic_vector(31 downto 0);
    signal NJ_265 : std_logic_vector(7 downto 0);
    signal NJ_265_251_buffered : std_logic_vector(7 downto 0);
    signal R_J_257_resized : std_logic_vector(7 downto 0);
    signal R_J_257_scaled : std_logic_vector(7 downto 0);
    signal ULT_u8_u1_269_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_258_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_258_final_offset : std_logic_vector(7 downto 0);
    signal array_obj_ref_258_offset_scale_factor_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_258_resized_base_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_258_root_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_258_word_address_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_258_word_offset_0 : std_logic_vector(7 downto 0);
    signal konst_263_wire_constant : std_logic_vector(7 downto 0);
    signal konst_268_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_250_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_258_offset_scale_factor_0 <= "00000001";
    array_obj_ref_258_resized_base_address <= "00000000";
    array_obj_ref_258_word_offset_0 <= "00000000";
    konst_263_wire_constant <= "00000001";
    konst_268_wire_constant <= "01000000";
    type_cast_250_wire_constant <= "00000000";
    phi_stmt_247: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_250_wire_constant & NJ_265_251_buffered;
      req <= phi_stmt_247_req_0 & phi_stmt_247_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_247",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_247_ack_0,
          idata => idata,
          odata => J_247,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_247
    NJ_265_251_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= NJ_265_251_buf_req_0;
      NJ_265_251_buf_ack_0<= wack(0);
      rreq(0) <= NJ_265_251_buf_req_1;
      NJ_265_251_buf_ack_1<= rack(0);
      NJ_265_251_buf : InterlockBuffer generic map ( -- 
        name => "NJ_265_251_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => NJ_265,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NJ_265_251_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_255_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_255_inst_req_0;
      type_cast_255_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_255_inst_req_1;
      type_cast_255_inst_ack_1<= rack(0);
      type_cast_255_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_255_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => J_247,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NJJ_256,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_258_addr_0
    process(array_obj_ref_258_root_address) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_258_root_address;
      ov(7 downto 0) := iv;
      array_obj_ref_258_word_address_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_258_gather_scatter
    process(NJJ_256) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := NJJ_256;
      ov(31 downto 0) := iv;
      array_obj_ref_258_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_258_index_0_rename
    process(R_J_257_resized) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_J_257_resized;
      ov(7 downto 0) := iv;
      R_J_257_scaled <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_258_index_0_resize
    process(J_247) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := J_247;
      ov(7 downto 0) := iv;
      R_J_257_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_258_index_offset
    process(R_J_257_scaled) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_J_257_scaled;
      ov(7 downto 0) := iv;
      array_obj_ref_258_final_offset <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_258_root_address_inst
    process(array_obj_ref_258_final_offset) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_258_final_offset;
      ov(7 downto 0) := iv;
      array_obj_ref_258_root_address <= ov(7 downto 0);
      --
    end process;
    if_stmt_266_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u8_u1_269_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_266_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_266_branch_req_0,
          ack0 => if_stmt_266_branch_ack_0,
          ack1 => if_stmt_266_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u8_u8_264_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= J_247;
      NJ_265 <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_264_inst_req_0;
      ADD_u8_u8_264_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_264_inst_req_1;
      ADD_u8_u8_264_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator ULT_u8_u1_269_inst
    process(J_247) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(J_247, konst_268_wire_constant, tmp_var);
      ULT_u8_u1_269_wire <= tmp_var; --
    end process;
    -- shared store operator group (0) : array_obj_ref_258_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(7 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_258_store_0_req_0;
      array_obj_ref_258_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_258_store_0_req_1;
      array_obj_ref_258_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_258_word_address_0;
      data_in <= array_obj_ref_258_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 8,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(7 downto 0),
          mdata => memory_space_2_sr_data(31 downto 0),
          mtag => memory_space_2_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end init_reg_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity jmp is -- 
  generic (tag_length : integer); 
  port ( -- 
    rs1_data : in  std_logic_vector(31 downto 0);
    pc : in  std_logic_vector(7 downto 0);
    next_pc : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity jmp;
architecture jmp_arch of jmp is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 40)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rs1_data_buffer :  std_logic_vector(31 downto 0);
  signal rs1_data_update_enable: Boolean;
  signal pc_buffer :  std_logic_vector(7 downto 0);
  signal pc_update_enable: Boolean;
  -- output port buffer signals
  signal next_pc_buffer :  std_logic_vector(7 downto 0);
  signal next_pc_update_enable: Boolean;
  signal jmp_CP_1177_start: Boolean;
  signal jmp_CP_1177_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal slice_280_inst_ack_1 : boolean;
  signal slice_280_inst_req_1 : boolean;
  signal slice_280_inst_req_0 : boolean;
  signal slice_280_inst_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "jmp_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 40) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= rs1_data;
  rs1_data_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(39 downto 32) <= pc;
  pc_buffer <= in_buffer_data_out(39 downto 32);
  in_buffer_data_in(tag_length + 39 downto 40) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 39 downto 40);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  jmp_CP_1177_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "jmp_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= next_pc_buffer;
  next_pc <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= jmp_CP_1177_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= jmp_CP_1177_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= jmp_CP_1177_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  jmp_CP_1177: Block -- control-path 
    signal jmp_CP_1177_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    jmp_CP_1177_elements(0) <= jmp_CP_1177_start;
    jmp_CP_1177_symbol <= jmp_CP_1177_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_281/slice_280_Update/$entry
      -- CP-element group 0: 	 assign_stmt_281/slice_280_Update/cr
      -- CP-element group 0: 	 assign_stmt_281/slice_280_Sample/rr
      -- CP-element group 0: 	 assign_stmt_281/slice_280_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_281/slice_280_update_start_
      -- CP-element group 0: 	 assign_stmt_281/slice_280_sample_start_
      -- CP-element group 0: 	 assign_stmt_281/$entry
      -- CP-element group 0: 	 $entry
      -- 
    rr_1190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => jmp_CP_1177_elements(0), ack => slice_280_inst_req_0); -- 
    cr_1195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => jmp_CP_1177_elements(0), ack => slice_280_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_281/slice_280_Sample/ra
      -- CP-element group 1: 	 assign_stmt_281/slice_280_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_281/slice_280_sample_completed_
      -- 
    ra_1191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_280_inst_ack_0, ack => jmp_CP_1177_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 assign_stmt_281/slice_280_Update/ca
      -- CP-element group 2: 	 assign_stmt_281/slice_280_Update/$exit
      -- CP-element group 2: 	 assign_stmt_281/slice_280_update_completed_
      -- CP-element group 2: 	 assign_stmt_281/$exit
      -- CP-element group 2: 	 $exit
      -- 
    ca_1196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_280_inst_ack_1, ack => jmp_CP_1177_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    -- 
  begin -- 
    slice_280_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_280_inst_req_0;
      slice_280_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_280_inst_req_1;
      slice_280_inst_ack_1<= update_ack(0);
      slice_280_inst: SliceSplitProtocol generic map(name => "slice_280_inst", in_data_width => 32, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => rs1_data_buffer, dout => next_pc_buffer, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- 
  end Block; -- data_path
  -- 
end jmp_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity load is -- 
  generic (tag_length : integer); 
  port ( -- 
    rs1_data : in  std_logic_vector(31 downto 0);
    rd : in  std_logic_vector(7 downto 0);
    pc : in  std_logic_vector(7 downto 0);
    next_pc : out  std_logic_vector(7 downto 0);
    accessMem_call_reqs : out  std_logic_vector(0 downto 0);
    accessMem_call_acks : in   std_logic_vector(0 downto 0);
    accessMem_call_data : out  std_logic_vector(40 downto 0);
    accessMem_call_tag  :  out  std_logic_vector(0 downto 0);
    accessMem_return_reqs : out  std_logic_vector(0 downto 0);
    accessMem_return_acks : in   std_logic_vector(0 downto 0);
    accessMem_return_data : in   std_logic_vector(31 downto 0);
    accessMem_return_tag :  in   std_logic_vector(0 downto 0);
    accessreg_call_reqs : out  std_logic_vector(0 downto 0);
    accessreg_call_acks : in   std_logic_vector(0 downto 0);
    accessreg_call_data : out  std_logic_vector(40 downto 0);
    accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
    accessreg_return_reqs : out  std_logic_vector(0 downto 0);
    accessreg_return_acks : in   std_logic_vector(0 downto 0);
    accessreg_return_data : in   std_logic_vector(31 downto 0);
    accessreg_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity load;
architecture load_arch of load is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 48)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rs1_data_buffer :  std_logic_vector(31 downto 0);
  signal rs1_data_update_enable: Boolean;
  signal rd_buffer :  std_logic_vector(7 downto 0);
  signal rd_update_enable: Boolean;
  signal pc_buffer :  std_logic_vector(7 downto 0);
  signal pc_update_enable: Boolean;
  -- output port buffer signals
  signal next_pc_buffer :  std_logic_vector(7 downto 0);
  signal next_pc_update_enable: Boolean;
  signal load_CP_1197_start: Boolean;
  signal load_CP_1197_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(7 downto 0);
      write_data : in  std_logic_vector(31 downto 0);
      read_data : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component accessreg is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(7 downto 0);
      write_data : in  std_logic_vector(31 downto 0);
      read_data : out  std_logic_vector(31 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_296_call_ack_0 : boolean;
  signal call_stmt_296_call_req_0 : boolean;
  signal call_stmt_301_call_req_0 : boolean;
  signal call_stmt_296_call_req_1 : boolean;
  signal call_stmt_296_call_ack_1 : boolean;
  signal ADD_u8_u8_305_inst_ack_1 : boolean;
  signal ADD_u8_u8_305_inst_req_1 : boolean;
  signal ADD_u8_u8_305_inst_ack_0 : boolean;
  signal ADD_u8_u8_305_inst_req_0 : boolean;
  signal call_stmt_301_call_ack_1 : boolean;
  signal call_stmt_301_call_req_1 : boolean;
  signal call_stmt_301_call_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "load_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 48) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= rs1_data;
  rs1_data_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(39 downto 32) <= rd;
  rd_buffer <= in_buffer_data_out(39 downto 32);
  in_buffer_data_in(47 downto 40) <= pc;
  pc_buffer <= in_buffer_data_out(47 downto 40);
  in_buffer_data_in(tag_length + 47 downto 48) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 47 downto 48);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  load_CP_1197_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "load_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= next_pc_buffer;
  next_pc <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= load_CP_1197_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= load_CP_1197_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= load_CP_1197_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  load_CP_1197: Block -- control-path 
    signal load_CP_1197_elements: BooleanArray(7 downto 0);
    -- 
  begin -- 
    load_CP_1197_elements(0) <= load_CP_1197_start;
    load_CP_1197_symbol <= load_CP_1197_elements(7);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0:  members (17) 
      -- CP-element group 0: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_301_update_start_
      -- CP-element group 0: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_296_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_296_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_296_sample_start_
      -- CP-element group 0: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_296_update_start_
      -- CP-element group 0: 	 assign_stmt_291_to_assign_stmt_306/$entry
      -- CP-element group 0: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_296_Sample/crr
      -- CP-element group 0: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_296_Update/ccr
      -- CP-element group 0: 	 assign_stmt_291_to_assign_stmt_306/ADD_u8_u8_305_Update/cr
      -- CP-element group 0: 	 assign_stmt_291_to_assign_stmt_306/ADD_u8_u8_305_Update/$entry
      -- CP-element group 0: 	 assign_stmt_291_to_assign_stmt_306/ADD_u8_u8_305_Sample/rr
      -- CP-element group 0: 	 assign_stmt_291_to_assign_stmt_306/ADD_u8_u8_305_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_291_to_assign_stmt_306/ADD_u8_u8_305_update_start_
      -- CP-element group 0: 	 assign_stmt_291_to_assign_stmt_306/ADD_u8_u8_305_sample_start_
      -- CP-element group 0: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_301_Update/ccr
      -- CP-element group 0: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_301_Update/$entry
      -- 
    crr_1210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => load_CP_1197_elements(0), ack => call_stmt_296_call_req_0); -- 
    ccr_1215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => load_CP_1197_elements(0), ack => call_stmt_296_call_req_1); -- 
    ccr_1229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => load_CP_1197_elements(0), ack => call_stmt_301_call_req_1); -- 
    rr_1238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => load_CP_1197_elements(0), ack => ADD_u8_u8_305_inst_req_0); -- 
    cr_1243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => load_CP_1197_elements(0), ack => ADD_u8_u8_305_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_296_Sample/cra
      -- CP-element group 1: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_296_sample_completed_
      -- CP-element group 1: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_296_Sample/$exit
      -- 
    cra_1211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_296_call_ack_0, ack => load_CP_1197_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_296_update_completed_
      -- CP-element group 2: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_296_Update/$exit
      -- CP-element group 2: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_301_Sample/crr
      -- CP-element group 2: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_296_Update/cca
      -- CP-element group 2: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_301_sample_start_
      -- CP-element group 2: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_301_Sample/$entry
      -- 
    cca_1216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_296_call_ack_1, ack => load_CP_1197_elements(2)); -- 
    crr_1224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => load_CP_1197_elements(2), ack => call_stmt_301_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_301_sample_completed_
      -- CP-element group 3: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_301_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_301_Sample/cra
      -- 
    cra_1225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_301_call_ack_0, ack => load_CP_1197_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_301_update_completed_
      -- CP-element group 4: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_301_Update/cca
      -- CP-element group 4: 	 assign_stmt_291_to_assign_stmt_306/call_stmt_301_Update/$exit
      -- 
    cca_1230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_301_call_ack_1, ack => load_CP_1197_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_291_to_assign_stmt_306/ADD_u8_u8_305_Sample/ra
      -- CP-element group 5: 	 assign_stmt_291_to_assign_stmt_306/ADD_u8_u8_305_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_291_to_assign_stmt_306/ADD_u8_u8_305_sample_completed_
      -- 
    ra_1239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_305_inst_ack_0, ack => load_CP_1197_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_291_to_assign_stmt_306/ADD_u8_u8_305_Update/ca
      -- CP-element group 6: 	 assign_stmt_291_to_assign_stmt_306/ADD_u8_u8_305_Update/$exit
      -- CP-element group 6: 	 assign_stmt_291_to_assign_stmt_306/ADD_u8_u8_305_update_completed_
      -- 
    ca_1244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_305_inst_ack_1, ack => load_CP_1197_elements(6)); -- 
    -- CP-element group 7:  join  transition  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 $exit
      -- CP-element group 7: 	 assign_stmt_291_to_assign_stmt_306/$exit
      -- 
    load_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 23) := "load_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= load_CP_1197_elements(4) & load_CP_1197_elements(6);
      gj_load_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => load_CP_1197_elements(7), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal addr_291 : std_logic_vector(7 downto 0);
    signal dummy1_301 : std_logic_vector(31 downto 0);
    signal konst_292_wire_constant : std_logic_vector(0 downto 0);
    signal konst_294_wire_constant : std_logic_vector(31 downto 0);
    signal konst_297_wire_constant : std_logic_vector(0 downto 0);
    signal konst_304_wire_constant : std_logic_vector(7 downto 0);
    signal output_296 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_292_wire_constant <= "1";
    konst_294_wire_constant <= "00000000000000000000000000000000";
    konst_297_wire_constant <= "0";
    konst_304_wire_constant <= "00000001";
    -- flow-through slice operator slice_290_inst
    addr_291 <= rs1_data_buffer(7 downto 0);
    -- shared split operator group (0) : ADD_u8_u8_305_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pc_buffer;
      next_pc_buffer <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_305_inst_req_0;
      ADD_u8_u8_305_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_305_inst_req_1;
      ADD_u8_u8_305_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared call operator group (0) : call_stmt_296_call 
    accessMem_call_group_0: Block -- 
      signal data_in: std_logic_vector(40 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_296_call_req_0;
      call_stmt_296_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_296_call_req_1;
      call_stmt_296_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMem_call_group_0_gI: SplitGuardInterface generic map(name => "accessMem_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_292_wire_constant & addr_291 & konst_294_wire_constant;
      output_296 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 41,
        owidth => 41,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMem_call_reqs(0),
          ackR => accessMem_call_acks(0),
          dataR => accessMem_call_data(40 downto 0),
          tagR => accessMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMem_return_acks(0), -- cross-over
          ackL => accessMem_return_reqs(0), -- cross-over
          dataL => accessMem_return_data(31 downto 0),
          tagL => accessMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_301_call 
    accessreg_call_group_1: Block -- 
      signal data_in: std_logic_vector(40 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_301_call_req_0;
      call_stmt_301_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_301_call_req_1;
      call_stmt_301_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessreg_call_group_1_gI: SplitGuardInterface generic map(name => "accessreg_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_297_wire_constant & rd_buffer & output_296;
      dummy1_301 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 41,
        owidth => 41,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessreg_call_reqs(0),
          ackR => accessreg_call_acks(0),
          dataR => accessreg_call_data(40 downto 0),
          tagR => accessreg_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessreg_return_acks(0), -- cross-over
          ackL => accessreg_return_reqs(0), -- cross-over
          dataL => accessreg_return_data(31 downto 0),
          tagL => accessreg_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end load_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity or_i is -- 
  generic (tag_length : integer); 
  port ( -- 
    rs1_data : in  std_logic_vector(31 downto 0);
    rs2_data : in  std_logic_vector(31 downto 0);
    rd : in  std_logic_vector(7 downto 0);
    pc : in  std_logic_vector(7 downto 0);
    next_pc : out  std_logic_vector(7 downto 0);
    accessreg_call_reqs : out  std_logic_vector(0 downto 0);
    accessreg_call_acks : in   std_logic_vector(0 downto 0);
    accessreg_call_data : out  std_logic_vector(40 downto 0);
    accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
    accessreg_return_reqs : out  std_logic_vector(0 downto 0);
    accessreg_return_acks : in   std_logic_vector(0 downto 0);
    accessreg_return_data : in   std_logic_vector(31 downto 0);
    accessreg_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity or_i;
architecture or_i_arch of or_i is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 80)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rs1_data_buffer :  std_logic_vector(31 downto 0);
  signal rs1_data_update_enable: Boolean;
  signal rs2_data_buffer :  std_logic_vector(31 downto 0);
  signal rs2_data_update_enable: Boolean;
  signal rd_buffer :  std_logic_vector(7 downto 0);
  signal rd_update_enable: Boolean;
  signal pc_buffer :  std_logic_vector(7 downto 0);
  signal pc_update_enable: Boolean;
  -- output port buffer signals
  signal next_pc_buffer :  std_logic_vector(7 downto 0);
  signal next_pc_update_enable: Boolean;
  signal or_i_CP_1245_start: Boolean;
  signal or_i_CP_1245_symbol: Boolean;
  -- volatile/operator module components. 
  component accessreg is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(7 downto 0);
      write_data : in  std_logic_vector(31 downto 0);
      read_data : out  std_logic_vector(31 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal ADD_u8_u8_327_inst_req_1 : boolean;
  signal ADD_u8_u8_327_inst_ack_1 : boolean;
  signal ADD_u8_u8_327_inst_req_0 : boolean;
  signal ADD_u8_u8_327_inst_ack_0 : boolean;
  signal call_stmt_323_call_ack_1 : boolean;
  signal call_stmt_323_call_req_1 : boolean;
  signal call_stmt_323_call_ack_0 : boolean;
  signal call_stmt_323_call_req_0 : boolean;
  signal OR_u32_u32_317_inst_ack_1 : boolean;
  signal OR_u32_u32_317_inst_req_1 : boolean;
  signal OR_u32_u32_317_inst_ack_0 : boolean;
  signal OR_u32_u32_317_inst_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "or_i_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 80) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= rs1_data;
  rs1_data_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= rs2_data;
  rs2_data_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(71 downto 64) <= rd;
  rd_buffer <= in_buffer_data_out(71 downto 64);
  in_buffer_data_in(79 downto 72) <= pc;
  pc_buffer <= in_buffer_data_out(79 downto 72);
  in_buffer_data_in(tag_length + 79 downto 80) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 79 downto 80);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  or_i_CP_1245_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "or_i_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= next_pc_buffer;
  next_pc <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= or_i_CP_1245_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= or_i_CP_1245_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= or_i_CP_1245_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  or_i_CP_1245: Block -- control-path 
    signal or_i_CP_1245_elements: BooleanArray(7 downto 0);
    -- 
  begin -- 
    or_i_CP_1245_elements(0) <= or_i_CP_1245_start;
    or_i_CP_1245_symbol <= or_i_CP_1245_elements(7);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0:  members (17) 
      -- CP-element group 0: 	 assign_stmt_318_to_assign_stmt_328/ADD_u8_u8_327_Update/cr
      -- CP-element group 0: 	 assign_stmt_318_to_assign_stmt_328/ADD_u8_u8_327_Update/$entry
      -- CP-element group 0: 	 assign_stmt_318_to_assign_stmt_328/ADD_u8_u8_327_Sample/rr
      -- CP-element group 0: 	 assign_stmt_318_to_assign_stmt_328/ADD_u8_u8_327_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_318_to_assign_stmt_328/ADD_u8_u8_327_update_start_
      -- CP-element group 0: 	 assign_stmt_318_to_assign_stmt_328/ADD_u8_u8_327_sample_start_
      -- CP-element group 0: 	 assign_stmt_318_to_assign_stmt_328/call_stmt_323_Update/ccr
      -- CP-element group 0: 	 assign_stmt_318_to_assign_stmt_328/call_stmt_323_Update/$entry
      -- CP-element group 0: 	 assign_stmt_318_to_assign_stmt_328/call_stmt_323_update_start_
      -- CP-element group 0: 	 assign_stmt_318_to_assign_stmt_328/OR_u32_u32_317_Update/cr
      -- CP-element group 0: 	 assign_stmt_318_to_assign_stmt_328/OR_u32_u32_317_Update/$entry
      -- CP-element group 0: 	 assign_stmt_318_to_assign_stmt_328/OR_u32_u32_317_Sample/rr
      -- CP-element group 0: 	 assign_stmt_318_to_assign_stmt_328/OR_u32_u32_317_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_318_to_assign_stmt_328/OR_u32_u32_317_update_start_
      -- CP-element group 0: 	 assign_stmt_318_to_assign_stmt_328/OR_u32_u32_317_sample_start_
      -- CP-element group 0: 	 assign_stmt_318_to_assign_stmt_328/$entry
      -- CP-element group 0: 	 $entry
      -- 
    rr_1258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => or_i_CP_1245_elements(0), ack => OR_u32_u32_317_inst_req_0); -- 
    cr_1263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => or_i_CP_1245_elements(0), ack => OR_u32_u32_317_inst_req_1); -- 
    ccr_1277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => or_i_CP_1245_elements(0), ack => call_stmt_323_call_req_1); -- 
    rr_1286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => or_i_CP_1245_elements(0), ack => ADD_u8_u8_327_inst_req_0); -- 
    cr_1291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => or_i_CP_1245_elements(0), ack => ADD_u8_u8_327_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_318_to_assign_stmt_328/OR_u32_u32_317_Sample/ra
      -- CP-element group 1: 	 assign_stmt_318_to_assign_stmt_328/OR_u32_u32_317_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_318_to_assign_stmt_328/OR_u32_u32_317_sample_completed_
      -- 
    ra_1259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_317_inst_ack_0, ack => or_i_CP_1245_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_318_to_assign_stmt_328/call_stmt_323_Sample/crr
      -- CP-element group 2: 	 assign_stmt_318_to_assign_stmt_328/call_stmt_323_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_318_to_assign_stmt_328/call_stmt_323_sample_start_
      -- CP-element group 2: 	 assign_stmt_318_to_assign_stmt_328/OR_u32_u32_317_Update/ca
      -- CP-element group 2: 	 assign_stmt_318_to_assign_stmt_328/OR_u32_u32_317_Update/$exit
      -- CP-element group 2: 	 assign_stmt_318_to_assign_stmt_328/OR_u32_u32_317_update_completed_
      -- 
    ca_1264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_317_inst_ack_1, ack => or_i_CP_1245_elements(2)); -- 
    crr_1272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => or_i_CP_1245_elements(2), ack => call_stmt_323_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_318_to_assign_stmt_328/call_stmt_323_Sample/cra
      -- CP-element group 3: 	 assign_stmt_318_to_assign_stmt_328/call_stmt_323_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_318_to_assign_stmt_328/call_stmt_323_sample_completed_
      -- 
    cra_1273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_323_call_ack_0, ack => or_i_CP_1245_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_318_to_assign_stmt_328/call_stmt_323_Update/cca
      -- CP-element group 4: 	 assign_stmt_318_to_assign_stmt_328/call_stmt_323_Update/$exit
      -- CP-element group 4: 	 assign_stmt_318_to_assign_stmt_328/call_stmt_323_update_completed_
      -- 
    cca_1278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_323_call_ack_1, ack => or_i_CP_1245_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_318_to_assign_stmt_328/ADD_u8_u8_327_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_318_to_assign_stmt_328/ADD_u8_u8_327_Sample/ra
      -- CP-element group 5: 	 assign_stmt_318_to_assign_stmt_328/ADD_u8_u8_327_sample_completed_
      -- 
    ra_1287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_327_inst_ack_0, ack => or_i_CP_1245_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_318_to_assign_stmt_328/ADD_u8_u8_327_Update/ca
      -- CP-element group 6: 	 assign_stmt_318_to_assign_stmt_328/ADD_u8_u8_327_Update/$exit
      -- CP-element group 6: 	 assign_stmt_318_to_assign_stmt_328/ADD_u8_u8_327_update_completed_
      -- 
    ca_1292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_327_inst_ack_1, ack => or_i_CP_1245_elements(6)); -- 
    -- CP-element group 7:  join  transition  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 assign_stmt_318_to_assign_stmt_328/$exit
      -- CP-element group 7: 	 $exit
      -- 
    or_i_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 23) := "or_i_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= or_i_CP_1245_elements(4) & or_i_CP_1245_elements(6);
      gj_or_i_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => or_i_CP_1245_elements(7), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal dummy_323 : std_logic_vector(31 downto 0);
    signal konst_319_wire_constant : std_logic_vector(0 downto 0);
    signal konst_326_wire_constant : std_logic_vector(7 downto 0);
    signal output_318 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_319_wire_constant <= "0";
    konst_326_wire_constant <= "00000001";
    -- shared split operator group (0) : ADD_u8_u8_327_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pc_buffer;
      next_pc_buffer <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_327_inst_req_0;
      ADD_u8_u8_327_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_327_inst_req_1;
      ADD_u8_u8_327_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : OR_u32_u32_317_inst 
    ApIntOr_group_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= rs1_data_buffer & rs2_data_buffer;
      output_318 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_317_inst_req_0;
      OR_u32_u32_317_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_317_inst_req_1;
      OR_u32_u32_317_inst_ack_1 <= ackR_unguarded(0);
      ApIntOr_group_1_gI: SplitGuardInterface generic map(name => "ApIntOr_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared call operator group (0) : call_stmt_323_call 
    accessreg_call_group_0: Block -- 
      signal data_in: std_logic_vector(40 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_323_call_req_0;
      call_stmt_323_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_323_call_req_1;
      call_stmt_323_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessreg_call_group_0_gI: SplitGuardInterface generic map(name => "accessreg_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_319_wire_constant & rd_buffer & output_318;
      dummy_323 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 41,
        owidth => 41,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessreg_call_reqs(0),
          ackR => accessreg_call_acks(0),
          dataR => accessreg_call_data(40 downto 0),
          tagR => accessreg_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessreg_return_acks(0), -- cross-over
          ackL => accessreg_return_reqs(0), -- cross-over
          dataL => accessreg_return_data(31 downto 0),
          tagL => accessreg_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end or_i_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sbir is -- 
  generic (tag_length : integer); 
  port ( -- 
    imm : in  std_logic_vector(7 downto 0);
    rd : in  std_logic_vector(7 downto 0);
    pc : in  std_logic_vector(7 downto 0);
    next_pc : out  std_logic_vector(7 downto 0);
    accessreg_call_reqs : out  std_logic_vector(0 downto 0);
    accessreg_call_acks : in   std_logic_vector(0 downto 0);
    accessreg_call_data : out  std_logic_vector(40 downto 0);
    accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
    accessreg_return_reqs : out  std_logic_vector(0 downto 0);
    accessreg_return_acks : in   std_logic_vector(0 downto 0);
    accessreg_return_data : in   std_logic_vector(31 downto 0);
    accessreg_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sbir;
architecture sbir_arch of sbir is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 24)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal imm_buffer :  std_logic_vector(7 downto 0);
  signal imm_update_enable: Boolean;
  signal rd_buffer :  std_logic_vector(7 downto 0);
  signal rd_update_enable: Boolean;
  signal pc_buffer :  std_logic_vector(7 downto 0);
  signal pc_update_enable: Boolean;
  -- output port buffer signals
  signal next_pc_buffer :  std_logic_vector(7 downto 0);
  signal next_pc_update_enable: Boolean;
  signal sbir_CP_1293_start: Boolean;
  signal sbir_CP_1293_symbol: Boolean;
  -- volatile/operator module components. 
  component accessreg is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(7 downto 0);
      write_data : in  std_logic_vector(31 downto 0);
      read_data : out  std_logic_vector(31 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_347_call_ack_0 : boolean;
  signal ADD_u8_u8_351_inst_ack_0 : boolean;
  signal call_stmt_347_call_req_0 : boolean;
  signal ADD_u8_u8_351_inst_req_1 : boolean;
  signal ADD_u8_u8_351_inst_ack_1 : boolean;
  signal CONCAT_u24_u32_341_inst_req_0 : boolean;
  signal CONCAT_u24_u32_341_inst_ack_0 : boolean;
  signal CONCAT_u24_u32_341_inst_req_1 : boolean;
  signal ADD_u8_u8_351_inst_req_0 : boolean;
  signal call_stmt_347_call_ack_1 : boolean;
  signal call_stmt_347_call_req_1 : boolean;
  signal CONCAT_u24_u32_341_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sbir_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 24) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= imm;
  imm_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(15 downto 8) <= rd;
  rd_buffer <= in_buffer_data_out(15 downto 8);
  in_buffer_data_in(23 downto 16) <= pc;
  pc_buffer <= in_buffer_data_out(23 downto 16);
  in_buffer_data_in(tag_length + 23 downto 24) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 23 downto 24);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sbir_CP_1293_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sbir_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= next_pc_buffer;
  next_pc <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sbir_CP_1293_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sbir_CP_1293_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sbir_CP_1293_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sbir_CP_1293: Block -- control-path 
    signal sbir_CP_1293_elements: BooleanArray(7 downto 0);
    -- 
  begin -- 
    sbir_CP_1293_elements(0) <= sbir_CP_1293_start;
    sbir_CP_1293_symbol <= sbir_CP_1293_elements(7);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0:  members (17) 
      -- CP-element group 0: 	 assign_stmt_342_to_assign_stmt_352/CONCAT_u24_u32_341_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_342_to_assign_stmt_352/$entry
      -- CP-element group 0: 	 assign_stmt_342_to_assign_stmt_352/CONCAT_u24_u32_341_sample_start_
      -- CP-element group 0: 	 assign_stmt_342_to_assign_stmt_352/call_stmt_347_update_start_
      -- CP-element group 0: 	 assign_stmt_342_to_assign_stmt_352/ADD_u8_u8_351_Update/$entry
      -- CP-element group 0: 	 assign_stmt_342_to_assign_stmt_352/call_stmt_347_Update/$entry
      -- CP-element group 0: 	 assign_stmt_342_to_assign_stmt_352/ADD_u8_u8_351_sample_start_
      -- CP-element group 0: 	 assign_stmt_342_to_assign_stmt_352/ADD_u8_u8_351_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_342_to_assign_stmt_352/ADD_u8_u8_351_Update/cr
      -- CP-element group 0: 	 assign_stmt_342_to_assign_stmt_352/CONCAT_u24_u32_341_Sample/rr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_342_to_assign_stmt_352/CONCAT_u24_u32_341_Update/$entry
      -- CP-element group 0: 	 assign_stmt_342_to_assign_stmt_352/CONCAT_u24_u32_341_Update/cr
      -- CP-element group 0: 	 assign_stmt_342_to_assign_stmt_352/ADD_u8_u8_351_Sample/rr
      -- CP-element group 0: 	 assign_stmt_342_to_assign_stmt_352/call_stmt_347_Update/ccr
      -- CP-element group 0: 	 assign_stmt_342_to_assign_stmt_352/ADD_u8_u8_351_update_start_
      -- CP-element group 0: 	 assign_stmt_342_to_assign_stmt_352/CONCAT_u24_u32_341_update_start_
      -- 
    rr_1306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sbir_CP_1293_elements(0), ack => CONCAT_u24_u32_341_inst_req_0); -- 
    cr_1311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sbir_CP_1293_elements(0), ack => CONCAT_u24_u32_341_inst_req_1); -- 
    ccr_1325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sbir_CP_1293_elements(0), ack => call_stmt_347_call_req_1); -- 
    rr_1334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sbir_CP_1293_elements(0), ack => ADD_u8_u8_351_inst_req_0); -- 
    cr_1339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sbir_CP_1293_elements(0), ack => ADD_u8_u8_351_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_342_to_assign_stmt_352/CONCAT_u24_u32_341_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_342_to_assign_stmt_352/CONCAT_u24_u32_341_Sample/ra
      -- CP-element group 1: 	 assign_stmt_342_to_assign_stmt_352/CONCAT_u24_u32_341_sample_completed_
      -- 
    ra_1307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u24_u32_341_inst_ack_0, ack => sbir_CP_1293_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_342_to_assign_stmt_352/CONCAT_u24_u32_341_update_completed_
      -- CP-element group 2: 	 assign_stmt_342_to_assign_stmt_352/call_stmt_347_sample_start_
      -- CP-element group 2: 	 assign_stmt_342_to_assign_stmt_352/CONCAT_u24_u32_341_Update/$exit
      -- CP-element group 2: 	 assign_stmt_342_to_assign_stmt_352/call_stmt_347_Sample/crr
      -- CP-element group 2: 	 assign_stmt_342_to_assign_stmt_352/call_stmt_347_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_342_to_assign_stmt_352/CONCAT_u24_u32_341_Update/ca
      -- 
    ca_1312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u24_u32_341_inst_ack_1, ack => sbir_CP_1293_elements(2)); -- 
    crr_1320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sbir_CP_1293_elements(2), ack => call_stmt_347_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_342_to_assign_stmt_352/call_stmt_347_Sample/cra
      -- CP-element group 3: 	 assign_stmt_342_to_assign_stmt_352/call_stmt_347_sample_completed_
      -- CP-element group 3: 	 assign_stmt_342_to_assign_stmt_352/call_stmt_347_Sample/$exit
      -- 
    cra_1321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_347_call_ack_0, ack => sbir_CP_1293_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_342_to_assign_stmt_352/call_stmt_347_update_completed_
      -- CP-element group 4: 	 assign_stmt_342_to_assign_stmt_352/call_stmt_347_Update/cca
      -- CP-element group 4: 	 assign_stmt_342_to_assign_stmt_352/call_stmt_347_Update/$exit
      -- 
    cca_1326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_347_call_ack_1, ack => sbir_CP_1293_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_342_to_assign_stmt_352/ADD_u8_u8_351_Sample/ra
      -- CP-element group 5: 	 assign_stmt_342_to_assign_stmt_352/ADD_u8_u8_351_sample_completed_
      -- CP-element group 5: 	 assign_stmt_342_to_assign_stmt_352/ADD_u8_u8_351_Sample/$exit
      -- 
    ra_1335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_351_inst_ack_0, ack => sbir_CP_1293_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_342_to_assign_stmt_352/ADD_u8_u8_351_update_completed_
      -- CP-element group 6: 	 assign_stmt_342_to_assign_stmt_352/ADD_u8_u8_351_Update/$exit
      -- CP-element group 6: 	 assign_stmt_342_to_assign_stmt_352/ADD_u8_u8_351_Update/ca
      -- 
    ca_1340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_351_inst_ack_1, ack => sbir_CP_1293_elements(6)); -- 
    -- CP-element group 7:  join  transition  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 assign_stmt_342_to_assign_stmt_352/$exit
      -- CP-element group 7: 	 $exit
      -- 
    sbir_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 23) := "sbir_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sbir_CP_1293_elements(4) & sbir_CP_1293_elements(6);
      gj_sbir_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sbir_CP_1293_elements(7), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_zero24_339_wire_constant : std_logic_vector(23 downto 0);
    signal dummy1_347 : std_logic_vector(31 downto 0);
    signal konst_343_wire_constant : std_logic_vector(0 downto 0);
    signal konst_350_wire_constant : std_logic_vector(7 downto 0);
    signal output_342 : std_logic_vector(31 downto 0);
    signal xxsbirxxzero24 : std_logic_vector(23 downto 0);
    -- 
  begin -- 
    R_zero24_339_wire_constant <= "000000000000000000000000";
    konst_343_wire_constant <= "0";
    konst_350_wire_constant <= "00000001";
    xxsbirxxzero24 <= "000000000000000000000000";
    -- shared split operator group (0) : ADD_u8_u8_351_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pc_buffer;
      next_pc_buffer <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_351_inst_req_0;
      ADD_u8_u8_351_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_351_inst_req_1;
      ADD_u8_u8_351_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : CONCAT_u24_u32_341_inst 
    ApConcat_group_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_zero24_339_wire_constant & imm_buffer;
      output_342 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u24_u32_341_inst_req_0;
      CONCAT_u24_u32_341_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u24_u32_341_inst_req_1;
      CONCAT_u24_u32_341_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_1_gI: SplitGuardInterface generic map(name => "ApConcat_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 24,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared call operator group (0) : call_stmt_347_call 
    accessreg_call_group_0: Block -- 
      signal data_in: std_logic_vector(40 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_347_call_req_0;
      call_stmt_347_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_347_call_req_1;
      call_stmt_347_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessreg_call_group_0_gI: SplitGuardInterface generic map(name => "accessreg_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_343_wire_constant & rd_buffer & output_342;
      dummy1_347 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 41,
        owidth => 41,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessreg_call_reqs(0),
          ackR => accessreg_call_acks(0),
          dataR => accessreg_call_data(40 downto 0),
          tagR => accessreg_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessreg_return_acks(0), -- cross-over
          ackL => accessreg_return_reqs(0), -- cross-over
          dataL => accessreg_return_data(31 downto 0),
          tagL => accessreg_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end sbir_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sll_i is -- 
  generic (tag_length : integer); 
  port ( -- 
    rs1_data : in  std_logic_vector(31 downto 0);
    rs2_data : in  std_logic_vector(31 downto 0);
    rd : in  std_logic_vector(7 downto 0);
    pc : in  std_logic_vector(7 downto 0);
    next_pc : out  std_logic_vector(7 downto 0);
    accessreg_call_reqs : out  std_logic_vector(0 downto 0);
    accessreg_call_acks : in   std_logic_vector(0 downto 0);
    accessreg_call_data : out  std_logic_vector(40 downto 0);
    accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
    accessreg_return_reqs : out  std_logic_vector(0 downto 0);
    accessreg_return_acks : in   std_logic_vector(0 downto 0);
    accessreg_return_data : in   std_logic_vector(31 downto 0);
    accessreg_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sll_i;
architecture sll_i_arch of sll_i is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 80)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rs1_data_buffer :  std_logic_vector(31 downto 0);
  signal rs1_data_update_enable: Boolean;
  signal rs2_data_buffer :  std_logic_vector(31 downto 0);
  signal rs2_data_update_enable: Boolean;
  signal rd_buffer :  std_logic_vector(7 downto 0);
  signal rd_update_enable: Boolean;
  signal pc_buffer :  std_logic_vector(7 downto 0);
  signal pc_update_enable: Boolean;
  -- output port buffer signals
  signal next_pc_buffer :  std_logic_vector(7 downto 0);
  signal next_pc_update_enable: Boolean;
  signal sll_i_CP_1341_start: Boolean;
  signal sll_i_CP_1341_symbol: Boolean;
  -- volatile/operator module components. 
  component accessreg is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(7 downto 0);
      write_data : in  std_logic_vector(31 downto 0);
      read_data : out  std_logic_vector(31 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal ADD_u8_u8_373_inst_ack_0 : boolean;
  signal ADD_u8_u8_373_inst_req_1 : boolean;
  signal call_stmt_369_call_ack_1 : boolean;
  signal ADD_u8_u8_373_inst_ack_1 : boolean;
  signal call_stmt_369_call_ack_0 : boolean;
  signal ADD_u8_u8_373_inst_req_0 : boolean;
  signal call_stmt_369_call_req_1 : boolean;
  signal call_stmt_369_call_req_0 : boolean;
  signal SHL_u32_u32_363_inst_ack_1 : boolean;
  signal SHL_u32_u32_363_inst_req_1 : boolean;
  signal SHL_u32_u32_363_inst_ack_0 : boolean;
  signal SHL_u32_u32_363_inst_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sll_i_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 80) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= rs1_data;
  rs1_data_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= rs2_data;
  rs2_data_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(71 downto 64) <= rd;
  rd_buffer <= in_buffer_data_out(71 downto 64);
  in_buffer_data_in(79 downto 72) <= pc;
  pc_buffer <= in_buffer_data_out(79 downto 72);
  in_buffer_data_in(tag_length + 79 downto 80) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 79 downto 80);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sll_i_CP_1341_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sll_i_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= next_pc_buffer;
  next_pc <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sll_i_CP_1341_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sll_i_CP_1341_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sll_i_CP_1341_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sll_i_CP_1341: Block -- control-path 
    signal sll_i_CP_1341_elements: BooleanArray(7 downto 0);
    -- 
  begin -- 
    sll_i_CP_1341_elements(0) <= sll_i_CP_1341_start;
    sll_i_CP_1341_symbol <= sll_i_CP_1341_elements(7);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0:  members (17) 
      -- CP-element group 0: 	 assign_stmt_364_to_assign_stmt_374/SHL_u32_u32_363_sample_start_
      -- CP-element group 0: 	 assign_stmt_364_to_assign_stmt_374/ADD_u8_u8_373_Update/cr
      -- CP-element group 0: 	 assign_stmt_364_to_assign_stmt_374/call_stmt_369_Update/$entry
      -- CP-element group 0: 	 assign_stmt_364_to_assign_stmt_374/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_364_to_assign_stmt_374/ADD_u8_u8_373_update_start_
      -- CP-element group 0: 	 assign_stmt_364_to_assign_stmt_374/SHL_u32_u32_363_update_start_
      -- CP-element group 0: 	 assign_stmt_364_to_assign_stmt_374/ADD_u8_u8_373_Sample/rr
      -- CP-element group 0: 	 assign_stmt_364_to_assign_stmt_374/ADD_u8_u8_373_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_364_to_assign_stmt_374/call_stmt_369_Update/ccr
      -- CP-element group 0: 	 assign_stmt_364_to_assign_stmt_374/ADD_u8_u8_373_Update/$entry
      -- CP-element group 0: 	 assign_stmt_364_to_assign_stmt_374/SHL_u32_u32_363_Update/cr
      -- CP-element group 0: 	 assign_stmt_364_to_assign_stmt_374/SHL_u32_u32_363_Update/$entry
      -- CP-element group 0: 	 assign_stmt_364_to_assign_stmt_374/SHL_u32_u32_363_Sample/rr
      -- CP-element group 0: 	 assign_stmt_364_to_assign_stmt_374/ADD_u8_u8_373_sample_start_
      -- CP-element group 0: 	 assign_stmt_364_to_assign_stmt_374/SHL_u32_u32_363_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_364_to_assign_stmt_374/call_stmt_369_update_start_
      -- 
    rr_1354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sll_i_CP_1341_elements(0), ack => SHL_u32_u32_363_inst_req_0); -- 
    cr_1359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sll_i_CP_1341_elements(0), ack => SHL_u32_u32_363_inst_req_1); -- 
    ccr_1373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sll_i_CP_1341_elements(0), ack => call_stmt_369_call_req_1); -- 
    rr_1382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sll_i_CP_1341_elements(0), ack => ADD_u8_u8_373_inst_req_0); -- 
    cr_1387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sll_i_CP_1341_elements(0), ack => ADD_u8_u8_373_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_364_to_assign_stmt_374/SHL_u32_u32_363_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_364_to_assign_stmt_374/SHL_u32_u32_363_sample_completed_
      -- CP-element group 1: 	 assign_stmt_364_to_assign_stmt_374/SHL_u32_u32_363_Sample/ra
      -- 
    ra_1355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_363_inst_ack_0, ack => sll_i_CP_1341_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_364_to_assign_stmt_374/call_stmt_369_sample_start_
      -- CP-element group 2: 	 assign_stmt_364_to_assign_stmt_374/SHL_u32_u32_363_update_completed_
      -- CP-element group 2: 	 assign_stmt_364_to_assign_stmt_374/call_stmt_369_Sample/crr
      -- CP-element group 2: 	 assign_stmt_364_to_assign_stmt_374/SHL_u32_u32_363_Update/ca
      -- CP-element group 2: 	 assign_stmt_364_to_assign_stmt_374/call_stmt_369_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_364_to_assign_stmt_374/SHL_u32_u32_363_Update/$exit
      -- 
    ca_1360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_363_inst_ack_1, ack => sll_i_CP_1341_elements(2)); -- 
    crr_1368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sll_i_CP_1341_elements(2), ack => call_stmt_369_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_364_to_assign_stmt_374/call_stmt_369_Sample/cra
      -- CP-element group 3: 	 assign_stmt_364_to_assign_stmt_374/call_stmt_369_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_364_to_assign_stmt_374/call_stmt_369_sample_completed_
      -- 
    cra_1369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_369_call_ack_0, ack => sll_i_CP_1341_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_364_to_assign_stmt_374/call_stmt_369_Update/cca
      -- CP-element group 4: 	 assign_stmt_364_to_assign_stmt_374/call_stmt_369_Update/$exit
      -- CP-element group 4: 	 assign_stmt_364_to_assign_stmt_374/call_stmt_369_update_completed_
      -- 
    cca_1374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_369_call_ack_1, ack => sll_i_CP_1341_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_364_to_assign_stmt_374/ADD_u8_u8_373_Sample/ra
      -- CP-element group 5: 	 assign_stmt_364_to_assign_stmt_374/ADD_u8_u8_373_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_364_to_assign_stmt_374/ADD_u8_u8_373_sample_completed_
      -- 
    ra_1383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_373_inst_ack_0, ack => sll_i_CP_1341_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_364_to_assign_stmt_374/ADD_u8_u8_373_Update/$exit
      -- CP-element group 6: 	 assign_stmt_364_to_assign_stmt_374/ADD_u8_u8_373_Update/ca
      -- CP-element group 6: 	 assign_stmt_364_to_assign_stmt_374/ADD_u8_u8_373_update_completed_
      -- 
    ca_1388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_373_inst_ack_1, ack => sll_i_CP_1341_elements(6)); -- 
    -- CP-element group 7:  join  transition  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 assign_stmt_364_to_assign_stmt_374/$exit
      -- CP-element group 7: 	 $exit
      -- 
    sll_i_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "sll_i_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sll_i_CP_1341_elements(4) & sll_i_CP_1341_elements(6);
      gj_sll_i_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sll_i_CP_1341_elements(7), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal dummy_369 : std_logic_vector(31 downto 0);
    signal konst_365_wire_constant : std_logic_vector(0 downto 0);
    signal konst_372_wire_constant : std_logic_vector(7 downto 0);
    signal output_364 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_365_wire_constant <= "0";
    konst_372_wire_constant <= "00000001";
    -- shared split operator group (0) : ADD_u8_u8_373_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pc_buffer;
      next_pc_buffer <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_373_inst_req_0;
      ADD_u8_u8_373_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_373_inst_req_1;
      ADD_u8_u8_373_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : SHL_u32_u32_363_inst 
    ApIntSHL_group_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= rs1_data_buffer & rs2_data_buffer;
      output_364 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SHL_u32_u32_363_inst_req_0;
      SHL_u32_u32_363_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_363_inst_req_1;
      SHL_u32_u32_363_inst_ack_1 <= ackR_unguarded(0);
      ApIntSHL_group_1_gI: SplitGuardInterface generic map(name => "ApIntSHL_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared call operator group (0) : call_stmt_369_call 
    accessreg_call_group_0: Block -- 
      signal data_in: std_logic_vector(40 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_369_call_req_0;
      call_stmt_369_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_369_call_req_1;
      call_stmt_369_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessreg_call_group_0_gI: SplitGuardInterface generic map(name => "accessreg_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_365_wire_constant & rd_buffer & output_364;
      dummy_369 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 41,
        owidth => 41,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessreg_call_reqs(0),
          ackR => accessreg_call_acks(0),
          dataR => accessreg_call_data(40 downto 0),
          tagR => accessreg_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessreg_return_acks(0), -- cross-over
          ackL => accessreg_return_reqs(0), -- cross-over
          dataL => accessreg_return_data(31 downto 0),
          tagL => accessreg_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end sll_i_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sra_i is -- 
  generic (tag_length : integer); 
  port ( -- 
    rs1_data : in  std_logic_vector(31 downto 0);
    rs2_data : in  std_logic_vector(31 downto 0);
    rd : in  std_logic_vector(7 downto 0);
    pc : in  std_logic_vector(7 downto 0);
    next_pc : out  std_logic_vector(7 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(2 downto 0);
    accessreg_call_reqs : out  std_logic_vector(0 downto 0);
    accessreg_call_acks : in   std_logic_vector(0 downto 0);
    accessreg_call_data : out  std_logic_vector(40 downto 0);
    accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
    accessreg_return_reqs : out  std_logic_vector(0 downto 0);
    accessreg_return_acks : in   std_logic_vector(0 downto 0);
    accessreg_return_data : in   std_logic_vector(31 downto 0);
    accessreg_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sra_i;
architecture sra_i_arch of sra_i is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 80)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rs1_data_buffer :  std_logic_vector(31 downto 0);
  signal rs1_data_update_enable: Boolean;
  signal rs2_data_buffer :  std_logic_vector(31 downto 0);
  signal rs2_data_update_enable: Boolean;
  signal rd_buffer :  std_logic_vector(7 downto 0);
  signal rd_update_enable: Boolean;
  signal pc_buffer :  std_logic_vector(7 downto 0);
  signal pc_update_enable: Boolean;
  -- output port buffer signals
  signal next_pc_buffer :  std_logic_vector(7 downto 0);
  signal next_pc_update_enable: Boolean;
  signal sra_i_CP_1389_start: Boolean;
  signal sra_i_CP_1389_symbol: Boolean;
  -- volatile/operator module components. 
  component accessreg is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(7 downto 0);
      write_data : in  std_logic_vector(31 downto 0);
      read_data : out  std_logic_vector(31 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal LSHR_u32_u32_385_inst_ack_0 : boolean;
  signal LSHR_u32_u32_385_inst_req_0 : boolean;
  signal LSHR_u32_u32_385_inst_req_1 : boolean;
  signal LSHR_u32_u32_385_inst_ack_1 : boolean;
  signal STORE_right_shift_382_store_0_req_0 : boolean;
  signal STORE_right_shift_382_store_0_ack_0 : boolean;
  signal STORE_right_shift_382_store_0_req_1 : boolean;
  signal STORE_right_shift_382_store_0_ack_1 : boolean;
  signal OR_u32_u32_400_inst_req_0 : boolean;
  signal OR_u32_u32_400_inst_ack_0 : boolean;
  signal OR_u32_u32_400_inst_req_1 : boolean;
  signal OR_u32_u32_400_inst_ack_1 : boolean;
  signal LOAD_right_shift_403_load_0_req_0 : boolean;
  signal LOAD_right_shift_403_load_0_ack_0 : boolean;
  signal LOAD_right_shift_403_load_0_req_1 : boolean;
  signal LOAD_right_shift_403_load_0_ack_1 : boolean;
  signal AND_u32_u32_405_inst_req_0 : boolean;
  signal AND_u32_u32_405_inst_ack_0 : boolean;
  signal AND_u32_u32_405_inst_req_1 : boolean;
  signal AND_u32_u32_405_inst_ack_1 : boolean;
  signal LOAD_right_shift_408_load_0_req_0 : boolean;
  signal LOAD_right_shift_408_load_0_ack_0 : boolean;
  signal LOAD_right_shift_408_load_0_req_1 : boolean;
  signal LOAD_right_shift_408_load_0_ack_1 : boolean;
  signal AND_u32_u32_411_inst_req_0 : boolean;
  signal AND_u32_u32_411_inst_ack_0 : boolean;
  signal AND_u32_u32_411_inst_req_1 : boolean;
  signal AND_u32_u32_411_inst_ack_1 : boolean;
  signal SHL_u32_u32_419_inst_req_0 : boolean;
  signal SHL_u32_u32_419_inst_ack_0 : boolean;
  signal SHL_u32_u32_419_inst_req_1 : boolean;
  signal SHL_u32_u32_419_inst_ack_1 : boolean;
  signal LOAD_right_shift_423_load_0_req_0 : boolean;
  signal LOAD_right_shift_423_load_0_ack_0 : boolean;
  signal LOAD_right_shift_423_load_0_req_1 : boolean;
  signal LOAD_right_shift_423_load_0_ack_1 : boolean;
  signal OR_u32_u32_425_inst_req_0 : boolean;
  signal OR_u32_u32_425_inst_ack_0 : boolean;
  signal OR_u32_u32_425_inst_req_1 : boolean;
  signal OR_u32_u32_425_inst_ack_1 : boolean;
  signal STORE_right_shift_422_store_0_req_0 : boolean;
  signal STORE_right_shift_422_store_0_ack_0 : boolean;
  signal STORE_right_shift_422_store_0_req_1 : boolean;
  signal STORE_right_shift_422_store_0_ack_1 : boolean;
  signal STORE_right_shift_428_store_0_req_0 : boolean;
  signal STORE_right_shift_428_store_0_ack_0 : boolean;
  signal STORE_right_shift_428_store_0_req_1 : boolean;
  signal STORE_right_shift_428_store_0_ack_1 : boolean;
  signal LOAD_right_shift_432_load_0_req_0 : boolean;
  signal LOAD_right_shift_432_load_0_ack_0 : boolean;
  signal LOAD_right_shift_432_load_0_req_1 : boolean;
  signal LOAD_right_shift_432_load_0_ack_1 : boolean;
  signal call_stmt_438_call_req_0 : boolean;
  signal call_stmt_438_call_ack_0 : boolean;
  signal call_stmt_438_call_req_1 : boolean;
  signal call_stmt_438_call_ack_1 : boolean;
  signal ADD_u8_u8_442_inst_req_0 : boolean;
  signal ADD_u8_u8_442_inst_ack_0 : boolean;
  signal ADD_u8_u8_442_inst_req_1 : boolean;
  signal ADD_u8_u8_442_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sra_i_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 80) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= rs1_data;
  rs1_data_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= rs2_data;
  rs2_data_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(71 downto 64) <= rd;
  rd_buffer <= in_buffer_data_out(71 downto 64);
  in_buffer_data_in(79 downto 72) <= pc;
  pc_buffer <= in_buffer_data_out(79 downto 72);
  in_buffer_data_in(tag_length + 79 downto 80) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 79 downto 80);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sra_i_CP_1389_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sra_i_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= next_pc_buffer;
  next_pc <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sra_i_CP_1389_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sra_i_CP_1389_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sra_i_CP_1389_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sra_i_CP_1389: Block -- control-path 
    signal sra_i_CP_1389_elements: BooleanArray(49 downto 0);
    -- 
  begin -- 
    sra_i_CP_1389_elements(0) <= sra_i_CP_1389_start;
    sra_i_CP_1389_symbol <= sra_i_CP_1389_elements(49);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	11 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	15 
    -- CP-element group 0: 	17 
    -- CP-element group 0: 	19 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	25 
    -- CP-element group 0: 	27 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	30 
    -- CP-element group 0: 	31 
    -- CP-element group 0: 	33 
    -- CP-element group 0: 	34 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	38 
    -- CP-element group 0: 	39 
    -- CP-element group 0: 	40 
    -- CP-element group 0:  members (84) 
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LSHR_u32_u32_385_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LSHR_u32_u32_385_Sample/rr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LSHR_u32_u32_385_update_start_
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LSHR_u32_u32_385_sample_start_
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LSHR_u32_u32_385_Update/cr
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_Update/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LSHR_u32_u32_385_Update/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_update_start_
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_400_sample_start_
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_400_update_start_
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_400_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_400_Sample/rr
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_400_Update/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_400_Update/cr
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_405_update_start_
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_update_start_
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_Update/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_405_Update/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_405_Update/cr
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_411_update_start_
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_update_start_
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_Update/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_411_Update/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_411_Update/cr
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/SHL_u32_u32_419_update_start_
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/SHL_u32_u32_419_Update/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/SHL_u32_u32_419_Update/cr
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_425_update_start_
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_update_start_
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_Update/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_425_Update/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_425_Update/cr
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_update_start_
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_Update/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_update_start_
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_Update/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_update_start_
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_Update/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/call_stmt_438_update_start_
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/call_stmt_438_Update/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/call_stmt_438_Update/ccr
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/ADD_u8_u8_442_sample_start_
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/ADD_u8_u8_442_update_start_
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/ADD_u8_u8_442_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/ADD_u8_u8_442_Sample/rr
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/ADD_u8_u8_442_Update/$entry
      -- CP-element group 0: 	 assign_stmt_386_to_assign_stmt_443/ADD_u8_u8_442_Update/cr
      -- 
    rr_1402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(0), ack => LSHR_u32_u32_385_inst_req_0); -- 
    cr_1407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(0), ack => LSHR_u32_u32_385_inst_req_1); -- 
    rr_1449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(0), ack => OR_u32_u32_400_inst_req_0); -- 
    cr_1454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(0), ack => OR_u32_u32_400_inst_req_1); -- 
    cr_1501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(0), ack => AND_u32_u32_405_inst_req_1); -- 
    cr_1486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(0), ack => LOAD_right_shift_403_load_0_req_1); -- 
    cr_1548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(0), ack => AND_u32_u32_411_inst_req_1); -- 
    cr_1533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(0), ack => LOAD_right_shift_408_load_0_req_1); -- 
    cr_1562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(0), ack => SHL_u32_u32_419_inst_req_1); -- 
    cr_1609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(0), ack => OR_u32_u32_425_inst_req_1); -- 
    cr_1594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(0), ack => LOAD_right_shift_423_load_0_req_1); -- 
    cr_1642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(0), ack => STORE_right_shift_422_store_0_req_1); -- 
    cr_1675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(0), ack => STORE_right_shift_428_store_0_req_1); -- 
    cr_1703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(0), ack => LOAD_right_shift_432_load_0_req_1); -- 
    ccr_1722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(0), ack => call_stmt_438_call_req_1); -- 
    rr_1731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(0), ack => ADD_u8_u8_442_inst_req_0); -- 
    cr_1736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(0), ack => ADD_u8_u8_442_inst_req_1); -- 
    cr_1440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(0), ack => STORE_right_shift_382_store_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_386_to_assign_stmt_443/LSHR_u32_u32_385_Sample/ra
      -- CP-element group 1: 	 assign_stmt_386_to_assign_stmt_443/LSHR_u32_u32_385_sample_completed_
      -- CP-element group 1: 	 assign_stmt_386_to_assign_stmt_443/LSHR_u32_u32_385_Sample/$exit
      -- 
    ra_1403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_385_inst_ack_0, ack => sra_i_CP_1389_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_386_to_assign_stmt_443/LSHR_u32_u32_385_update_completed_
      -- CP-element group 2: 	 assign_stmt_386_to_assign_stmt_443/LSHR_u32_u32_385_Update/ca
      -- CP-element group 2: 	 assign_stmt_386_to_assign_stmt_443/LSHR_u32_u32_385_Update/$exit
      -- 
    ca_1408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_385_inst_ack_1, ack => sra_i_CP_1389_elements(2)); -- 
    -- CP-element group 3:  join  transition  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_sample_start_
      -- CP-element group 3: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_Sample/$entry
      -- CP-element group 3: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_Sample/STORE_right_shift_382_Split/$entry
      -- CP-element group 3: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_Sample/STORE_right_shift_382_Split/$exit
      -- CP-element group 3: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_Sample/word_access_start/word_0/rr
      -- CP-element group 3: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_Sample/word_access_start/$entry
      -- CP-element group 3: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_Sample/STORE_right_shift_382_Split/split_req
      -- CP-element group 3: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_Sample/STORE_right_shift_382_Split/split_ack
      -- 
    rr_1429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(3), ack => STORE_right_shift_382_store_0_req_0); -- 
    sra_i_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "sra_i_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sra_i_CP_1389_elements(0) & sra_i_CP_1389_elements(2);
      gj_sra_i_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sra_i_CP_1389_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  fork  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	41 
    -- CP-element group 4: 	42 
    -- CP-element group 4: 	43 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_Sample/$exit
      -- CP-element group 4: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_Sample/word_access_start/word_0/ra
      -- CP-element group 4: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_Sample/word_access_start/$exit
      -- CP-element group 4: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_Sample/word_access_start/word_0/$exit
      -- CP-element group 4: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_sample_completed_
      -- 
    ra_1430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_right_shift_382_store_0_ack_0, ack => sra_i_CP_1389_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	49 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_Update/$exit
      -- CP-element group 5: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_Update/word_access_complete/$exit
      -- CP-element group 5: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_update_completed_
      -- CP-element group 5: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_Update/word_access_complete/word_0/$exit
      -- CP-element group 5: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_Update/word_access_complete/word_0/ca
      -- 
    ca_1441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_right_shift_382_store_0_ack_1, ack => sra_i_CP_1389_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_400_sample_completed_
      -- CP-element group 6: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_400_Sample/$exit
      -- CP-element group 6: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_400_Sample/ra
      -- 
    ra_1450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_400_inst_ack_0, ack => sra_i_CP_1389_elements(6)); -- 
    -- CP-element group 7:  fork  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7: 	14 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_400_update_completed_
      -- CP-element group 7: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_400_Update/$exit
      -- CP-element group 7: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_400_Update/ca
      -- 
    ca_1455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_400_inst_ack_1, ack => sra_i_CP_1389_elements(7)); -- 
    -- CP-element group 8:  join  transition  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: 	11 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	12 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_405_sample_start_
      -- CP-element group 8: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_405_Sample/$entry
      -- CP-element group 8: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_405_Sample/rr
      -- 
    rr_1496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(8), ack => AND_u32_u32_405_inst_req_0); -- 
    sra_i_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "sra_i_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sra_i_CP_1389_elements(7) & sra_i_CP_1389_elements(11);
      gj_sra_i_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sra_i_CP_1389_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  transition  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: 	41 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_sample_start_
      -- CP-element group 9: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_Sample/$entry
      -- CP-element group 9: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_Sample/word_access_start/$entry
      -- CP-element group 9: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_Sample/word_access_start/word_0/$entry
      -- CP-element group 9: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_Sample/word_access_start/word_0/rr
      -- 
    rr_1475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(9), ack => LOAD_right_shift_403_load_0_req_0); -- 
    sra_i_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "sra_i_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sra_i_CP_1389_elements(0) & sra_i_CP_1389_elements(41);
      gj_sra_i_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sra_i_CP_1389_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	44 
    -- CP-element group 10:  members (5) 
      -- CP-element group 10: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_sample_completed_
      -- CP-element group 10: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_Sample/$exit
      -- CP-element group 10: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_Sample/word_access_start/$exit
      -- CP-element group 10: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_Sample/word_access_start/word_0/$exit
      -- CP-element group 10: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_Sample/word_access_start/word_0/ra
      -- 
    ra_1476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_right_shift_403_load_0_ack_0, ack => sra_i_CP_1389_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	8 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_update_completed_
      -- CP-element group 11: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_Update/$exit
      -- CP-element group 11: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_Update/word_access_complete/$exit
      -- CP-element group 11: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_Update/word_access_complete/word_0/$exit
      -- CP-element group 11: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_Update/word_access_complete/word_0/ca
      -- CP-element group 11: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_Update/LOAD_right_shift_403_Merge/$entry
      -- CP-element group 11: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_Update/LOAD_right_shift_403_Merge/$exit
      -- CP-element group 11: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_Update/LOAD_right_shift_403_Merge/merge_req
      -- CP-element group 11: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_Update/LOAD_right_shift_403_Merge/merge_ack
      -- 
    ca_1487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_right_shift_403_load_0_ack_1, ack => sra_i_CP_1389_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	8 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_405_sample_completed_
      -- CP-element group 12: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_405_Sample/$exit
      -- CP-element group 12: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_405_Sample/ra
      -- 
    ra_1497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_405_inst_ack_0, ack => sra_i_CP_1389_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	20 
    -- CP-element group 13: 	22 
    -- CP-element group 13: 	23 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_405_update_completed_
      -- CP-element group 13: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_405_Update/$exit
      -- CP-element group 13: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_405_Update/ca
      -- CP-element group 13: 	 assign_stmt_386_to_assign_stmt_443/SHL_u32_u32_419_sample_start_
      -- CP-element group 13: 	 assign_stmt_386_to_assign_stmt_443/SHL_u32_u32_419_Sample/$entry
      -- CP-element group 13: 	 assign_stmt_386_to_assign_stmt_443/SHL_u32_u32_419_Sample/rr
      -- 
    ca_1502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_405_inst_ack_1, ack => sra_i_CP_1389_elements(13)); -- 
    rr_1557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(13), ack => SHL_u32_u32_419_inst_req_0); -- 
    -- CP-element group 14:  join  transition  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	7 
    -- CP-element group 14: 	17 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	18 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_411_sample_start_
      -- CP-element group 14: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_411_Sample/$entry
      -- CP-element group 14: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_411_Sample/rr
      -- 
    rr_1543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(14), ack => AND_u32_u32_411_inst_req_0); -- 
    sra_i_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sra_i_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sra_i_CP_1389_elements(7) & sra_i_CP_1389_elements(17);
      gj_sra_i_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sra_i_CP_1389_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	0 
    -- CP-element group 15: 	42 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_sample_start_
      -- CP-element group 15: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_Sample/$entry
      -- CP-element group 15: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_Sample/word_access_start/$entry
      -- CP-element group 15: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_Sample/word_access_start/word_0/$entry
      -- CP-element group 15: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_Sample/word_access_start/word_0/rr
      -- 
    rr_1522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(15), ack => LOAD_right_shift_408_load_0_req_0); -- 
    sra_i_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sra_i_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sra_i_CP_1389_elements(0) & sra_i_CP_1389_elements(42);
      gj_sra_i_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sra_i_CP_1389_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	45 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_sample_completed_
      -- CP-element group 16: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_Sample/$exit
      -- CP-element group 16: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_Sample/word_access_start/$exit
      -- CP-element group 16: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_Sample/word_access_start/word_0/$exit
      -- CP-element group 16: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_Sample/word_access_start/word_0/ra
      -- 
    ra_1523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_right_shift_408_load_0_ack_0, ack => sra_i_CP_1389_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	14 
    -- CP-element group 17:  members (9) 
      -- CP-element group 17: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_update_completed_
      -- CP-element group 17: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_Update/$exit
      -- CP-element group 17: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_Update/word_access_complete/$exit
      -- CP-element group 17: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_Update/word_access_complete/word_0/$exit
      -- CP-element group 17: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_Update/word_access_complete/word_0/ca
      -- CP-element group 17: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_Update/LOAD_right_shift_408_Merge/$entry
      -- CP-element group 17: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_Update/LOAD_right_shift_408_Merge/$exit
      -- CP-element group 17: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_Update/LOAD_right_shift_408_Merge/merge_req
      -- CP-element group 17: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_Update/LOAD_right_shift_408_Merge/merge_ack
      -- 
    ca_1534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_right_shift_408_load_0_ack_1, ack => sra_i_CP_1389_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_411_sample_completed_
      -- CP-element group 18: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_411_Sample/$exit
      -- CP-element group 18: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_411_Sample/ra
      -- 
    ra_1544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_411_inst_ack_0, ack => sra_i_CP_1389_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	0 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	31 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_411_update_completed_
      -- CP-element group 19: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_411_Update/$exit
      -- CP-element group 19: 	 assign_stmt_386_to_assign_stmt_443/AND_u32_u32_411_Update/ca
      -- 
    ca_1549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u32_u32_411_inst_ack_1, ack => sra_i_CP_1389_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	13 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 assign_stmt_386_to_assign_stmt_443/SHL_u32_u32_419_sample_completed_
      -- CP-element group 20: 	 assign_stmt_386_to_assign_stmt_443/SHL_u32_u32_419_Sample/$exit
      -- CP-element group 20: 	 assign_stmt_386_to_assign_stmt_443/SHL_u32_u32_419_Sample/ra
      -- 
    ra_1558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_419_inst_ack_0, ack => sra_i_CP_1389_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 assign_stmt_386_to_assign_stmt_443/SHL_u32_u32_419_update_completed_
      -- CP-element group 21: 	 assign_stmt_386_to_assign_stmt_443/SHL_u32_u32_419_Update/$exit
      -- CP-element group 21: 	 assign_stmt_386_to_assign_stmt_443/SHL_u32_u32_419_Update/ca
      -- 
    ca_1563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SHL_u32_u32_419_inst_ack_1, ack => sra_i_CP_1389_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	13 
    -- CP-element group 22: 	21 
    -- CP-element group 22: 	25 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	26 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_425_sample_start_
      -- CP-element group 22: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_425_Sample/$entry
      -- CP-element group 22: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_425_Sample/rr
      -- 
    rr_1604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(22), ack => OR_u32_u32_425_inst_req_0); -- 
    sra_i_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sra_i_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sra_i_CP_1389_elements(13) & sra_i_CP_1389_elements(21) & sra_i_CP_1389_elements(25);
      gj_sra_i_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sra_i_CP_1389_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: 	13 
    -- CP-element group 23: 	43 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_sample_start_
      -- CP-element group 23: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_Sample/$entry
      -- CP-element group 23: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_Sample/word_access_start/$entry
      -- CP-element group 23: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_Sample/word_access_start/word_0/$entry
      -- CP-element group 23: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_Sample/word_access_start/word_0/rr
      -- 
    rr_1583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(23), ack => LOAD_right_shift_423_load_0_req_0); -- 
    sra_i_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sra_i_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sra_i_CP_1389_elements(0) & sra_i_CP_1389_elements(13) & sra_i_CP_1389_elements(43);
      gj_sra_i_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sra_i_CP_1389_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	46 
    -- CP-element group 24:  members (5) 
      -- CP-element group 24: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_sample_completed_
      -- CP-element group 24: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_Sample/$exit
      -- CP-element group 24: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_Sample/word_access_start/$exit
      -- CP-element group 24: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_Sample/word_access_start/word_0/$exit
      -- CP-element group 24: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_Sample/word_access_start/word_0/ra
      -- 
    ra_1584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_right_shift_423_load_0_ack_0, ack => sra_i_CP_1389_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	0 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	22 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_update_completed_
      -- CP-element group 25: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_Update/$exit
      -- CP-element group 25: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_Update/word_access_complete/$exit
      -- CP-element group 25: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_Update/word_access_complete/word_0/$exit
      -- CP-element group 25: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_Update/word_access_complete/word_0/ca
      -- CP-element group 25: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_Update/LOAD_right_shift_423_Merge/$entry
      -- CP-element group 25: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_Update/LOAD_right_shift_423_Merge/$exit
      -- CP-element group 25: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_Update/LOAD_right_shift_423_Merge/merge_req
      -- CP-element group 25: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_Update/LOAD_right_shift_423_Merge/merge_ack
      -- 
    ca_1595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_right_shift_423_load_0_ack_1, ack => sra_i_CP_1389_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	22 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_425_sample_completed_
      -- CP-element group 26: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_425_Sample/$exit
      -- CP-element group 26: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_425_Sample/ra
      -- 
    ra_1605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_425_inst_ack_0, ack => sra_i_CP_1389_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_425_update_completed_
      -- CP-element group 27: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_425_Update/$exit
      -- CP-element group 27: 	 assign_stmt_386_to_assign_stmt_443/OR_u32_u32_425_Update/ca
      -- 
    ca_1610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u32_u32_425_inst_ack_1, ack => sra_i_CP_1389_elements(27)); -- 
    -- CP-element group 28:  join  transition  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: 	27 
    -- CP-element group 28: 	44 
    -- CP-element group 28: 	45 
    -- CP-element group 28: 	46 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_sample_start_
      -- CP-element group 28: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_Sample/$entry
      -- CP-element group 28: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_Sample/STORE_right_shift_422_Split/$entry
      -- CP-element group 28: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_Sample/STORE_right_shift_422_Split/$exit
      -- CP-element group 28: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_Sample/STORE_right_shift_422_Split/split_req
      -- CP-element group 28: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_Sample/STORE_right_shift_422_Split/split_ack
      -- CP-element group 28: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_Sample/word_access_start/$entry
      -- CP-element group 28: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_Sample/word_access_start/word_0/$entry
      -- CP-element group 28: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_Sample/word_access_start/word_0/rr
      -- 
    rr_1631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(28), ack => STORE_right_shift_422_store_0_req_0); -- 
    sra_i_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 25) := "sra_i_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= sra_i_CP_1389_elements(0) & sra_i_CP_1389_elements(27) & sra_i_CP_1389_elements(44) & sra_i_CP_1389_elements(45) & sra_i_CP_1389_elements(46);
      gj_sra_i_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sra_i_CP_1389_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	47 
    -- CP-element group 29:  members (5) 
      -- CP-element group 29: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_sample_completed_
      -- CP-element group 29: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_Sample/$exit
      -- CP-element group 29: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_Sample/word_access_start/$exit
      -- CP-element group 29: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_Sample/word_access_start/word_0/$exit
      -- CP-element group 29: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_Sample/word_access_start/word_0/ra
      -- 
    ra_1632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_right_shift_422_store_0_ack_0, ack => sra_i_CP_1389_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	0 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	49 
    -- CP-element group 30:  members (5) 
      -- CP-element group 30: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_update_completed_
      -- CP-element group 30: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_Update/$exit
      -- CP-element group 30: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_Update/word_access_complete/$exit
      -- CP-element group 30: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_Update/word_access_complete/word_0/$exit
      -- CP-element group 30: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_Update/word_access_complete/word_0/ca
      -- 
    ca_1643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_right_shift_422_store_0_ack_1, ack => sra_i_CP_1389_elements(30)); -- 
    -- CP-element group 31:  join  transition  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	0 
    -- CP-element group 31: 	19 
    -- CP-element group 31: 	47 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_sample_start_
      -- CP-element group 31: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_Sample/$entry
      -- CP-element group 31: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_Sample/STORE_right_shift_428_Split/$entry
      -- CP-element group 31: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_Sample/STORE_right_shift_428_Split/$exit
      -- CP-element group 31: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_Sample/STORE_right_shift_428_Split/split_req
      -- CP-element group 31: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_Sample/STORE_right_shift_428_Split/split_ack
      -- CP-element group 31: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_Sample/word_access_start/$entry
      -- CP-element group 31: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_Sample/word_access_start/word_0/$entry
      -- CP-element group 31: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_Sample/word_access_start/word_0/rr
      -- 
    rr_1664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(31), ack => STORE_right_shift_428_store_0_req_0); -- 
    sra_i_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sra_i_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sra_i_CP_1389_elements(0) & sra_i_CP_1389_elements(19) & sra_i_CP_1389_elements(47);
      gj_sra_i_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sra_i_CP_1389_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	48 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_sample_completed_
      -- CP-element group 32: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_Sample/$exit
      -- CP-element group 32: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_Sample/word_access_start/$exit
      -- CP-element group 32: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_Sample/word_access_start/word_0/$exit
      -- CP-element group 32: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_Sample/word_access_start/word_0/ra
      -- 
    ra_1665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_right_shift_428_store_0_ack_0, ack => sra_i_CP_1389_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	0 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	49 
    -- CP-element group 33:  members (5) 
      -- CP-element group 33: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_update_completed_
      -- CP-element group 33: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_Update/$exit
      -- CP-element group 33: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_Update/word_access_complete/$exit
      -- CP-element group 33: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_Update/word_access_complete/word_0/$exit
      -- CP-element group 33: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_Update/word_access_complete/word_0/ca
      -- 
    ca_1676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_right_shift_428_store_0_ack_1, ack => sra_i_CP_1389_elements(33)); -- 
    -- CP-element group 34:  join  transition  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	0 
    -- CP-element group 34: 	48 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_sample_start_
      -- CP-element group 34: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_Sample/$entry
      -- CP-element group 34: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_Sample/word_access_start/$entry
      -- CP-element group 34: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_Sample/word_access_start/word_0/$entry
      -- CP-element group 34: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_Sample/word_access_start/word_0/rr
      -- 
    rr_1692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(34), ack => LOAD_right_shift_432_load_0_req_0); -- 
    sra_i_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sra_i_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sra_i_CP_1389_elements(0) & sra_i_CP_1389_elements(48);
      gj_sra_i_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sra_i_CP_1389_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (5) 
      -- CP-element group 35: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_sample_completed_
      -- CP-element group 35: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_Sample/$exit
      -- CP-element group 35: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_Sample/word_access_start/$exit
      -- CP-element group 35: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_Sample/word_access_start/word_0/$exit
      -- CP-element group 35: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_Sample/word_access_start/word_0/ra
      -- 
    ra_1693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_right_shift_432_load_0_ack_0, ack => sra_i_CP_1389_elements(35)); -- 
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (12) 
      -- CP-element group 36: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_update_completed_
      -- CP-element group 36: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_Update/$exit
      -- CP-element group 36: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_Update/word_access_complete/$exit
      -- CP-element group 36: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_Update/word_access_complete/word_0/$exit
      -- CP-element group 36: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_Update/word_access_complete/word_0/ca
      -- CP-element group 36: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_Update/LOAD_right_shift_432_Merge/$entry
      -- CP-element group 36: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_Update/LOAD_right_shift_432_Merge/$exit
      -- CP-element group 36: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_Update/LOAD_right_shift_432_Merge/merge_req
      -- CP-element group 36: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_432_Update/LOAD_right_shift_432_Merge/merge_ack
      -- CP-element group 36: 	 assign_stmt_386_to_assign_stmt_443/call_stmt_438_sample_start_
      -- CP-element group 36: 	 assign_stmt_386_to_assign_stmt_443/call_stmt_438_Sample/$entry
      -- CP-element group 36: 	 assign_stmt_386_to_assign_stmt_443/call_stmt_438_Sample/crr
      -- 
    ca_1704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_right_shift_432_load_0_ack_1, ack => sra_i_CP_1389_elements(36)); -- 
    crr_1717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sra_i_CP_1389_elements(36), ack => call_stmt_438_call_req_0); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 assign_stmt_386_to_assign_stmt_443/call_stmt_438_sample_completed_
      -- CP-element group 37: 	 assign_stmt_386_to_assign_stmt_443/call_stmt_438_Sample/$exit
      -- CP-element group 37: 	 assign_stmt_386_to_assign_stmt_443/call_stmt_438_Sample/cra
      -- 
    cra_1718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_438_call_ack_0, ack => sra_i_CP_1389_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	0 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	49 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 assign_stmt_386_to_assign_stmt_443/call_stmt_438_update_completed_
      -- CP-element group 38: 	 assign_stmt_386_to_assign_stmt_443/call_stmt_438_Update/$exit
      -- CP-element group 38: 	 assign_stmt_386_to_assign_stmt_443/call_stmt_438_Update/cca
      -- 
    cca_1723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_438_call_ack_1, ack => sra_i_CP_1389_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	0 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 assign_stmt_386_to_assign_stmt_443/ADD_u8_u8_442_sample_completed_
      -- CP-element group 39: 	 assign_stmt_386_to_assign_stmt_443/ADD_u8_u8_442_Sample/$exit
      -- CP-element group 39: 	 assign_stmt_386_to_assign_stmt_443/ADD_u8_u8_442_Sample/ra
      -- 
    ra_1732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_442_inst_ack_0, ack => sra_i_CP_1389_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	49 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 assign_stmt_386_to_assign_stmt_443/ADD_u8_u8_442_update_completed_
      -- CP-element group 40: 	 assign_stmt_386_to_assign_stmt_443/ADD_u8_u8_442_Update/$exit
      -- CP-element group 40: 	 assign_stmt_386_to_assign_stmt_443/ADD_u8_u8_442_Update/ca
      -- 
    ca_1737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_442_inst_ack_1, ack => sra_i_CP_1389_elements(40)); -- 
    -- CP-element group 41:  transition  delay-element  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	4 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	9 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_LOAD_right_shift_403_delay
      -- 
    -- Element group sra_i_CP_1389_elements(41) is a control-delay.
    cp_element_41_delay: control_delay_element  generic map(name => " 41_delay", delay_value => 1)  port map(req => sra_i_CP_1389_elements(4), ack => sra_i_CP_1389_elements(41), clk => clk, reset =>reset);
    -- CP-element group 42:  transition  delay-element  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	4 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	15 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_LOAD_right_shift_408_delay
      -- 
    -- Element group sra_i_CP_1389_elements(42) is a control-delay.
    cp_element_42_delay: control_delay_element  generic map(name => " 42_delay", delay_value => 1)  port map(req => sra_i_CP_1389_elements(4), ack => sra_i_CP_1389_elements(42), clk => clk, reset =>reset);
    -- CP-element group 43:  transition  delay-element  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	4 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	23 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_382_LOAD_right_shift_423_delay
      -- 
    -- Element group sra_i_CP_1389_elements(43) is a control-delay.
    cp_element_43_delay: control_delay_element  generic map(name => " 43_delay", delay_value => 1)  port map(req => sra_i_CP_1389_elements(4), ack => sra_i_CP_1389_elements(43), clk => clk, reset =>reset);
    -- CP-element group 44:  transition  delay-element  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	10 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	28 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_403_STORE_right_shift_422_delay
      -- 
    -- Element group sra_i_CP_1389_elements(44) is a control-delay.
    cp_element_44_delay: control_delay_element  generic map(name => " 44_delay", delay_value => 1)  port map(req => sra_i_CP_1389_elements(10), ack => sra_i_CP_1389_elements(44), clk => clk, reset =>reset);
    -- CP-element group 45:  transition  delay-element  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	16 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	28 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_408_STORE_right_shift_422_delay
      -- 
    -- Element group sra_i_CP_1389_elements(45) is a control-delay.
    cp_element_45_delay: control_delay_element  generic map(name => " 45_delay", delay_value => 1)  port map(req => sra_i_CP_1389_elements(16), ack => sra_i_CP_1389_elements(45), clk => clk, reset =>reset);
    -- CP-element group 46:  transition  delay-element  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	24 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	28 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 assign_stmt_386_to_assign_stmt_443/LOAD_right_shift_423_STORE_right_shift_422_delay
      -- 
    -- Element group sra_i_CP_1389_elements(46) is a control-delay.
    cp_element_46_delay: control_delay_element  generic map(name => " 46_delay", delay_value => 1)  port map(req => sra_i_CP_1389_elements(24), ack => sra_i_CP_1389_elements(46), clk => clk, reset =>reset);
    -- CP-element group 47:  transition  delay-element  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	29 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	31 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_422_STORE_right_shift_428_delay
      -- 
    -- Element group sra_i_CP_1389_elements(47) is a control-delay.
    cp_element_47_delay: control_delay_element  generic map(name => " 47_delay", delay_value => 1)  port map(req => sra_i_CP_1389_elements(29), ack => sra_i_CP_1389_elements(47), clk => clk, reset =>reset);
    -- CP-element group 48:  transition  delay-element  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	32 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	34 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 assign_stmt_386_to_assign_stmt_443/STORE_right_shift_428_LOAD_right_shift_432_delay
      -- 
    -- Element group sra_i_CP_1389_elements(48) is a control-delay.
    cp_element_48_delay: control_delay_element  generic map(name => " 48_delay", delay_value => 1)  port map(req => sra_i_CP_1389_elements(32), ack => sra_i_CP_1389_elements(48), clk => clk, reset =>reset);
    -- CP-element group 49:  join  transition  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	5 
    -- CP-element group 49: 	30 
    -- CP-element group 49: 	33 
    -- CP-element group 49: 	38 
    -- CP-element group 49: 	40 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 assign_stmt_386_to_assign_stmt_443/$exit
      -- CP-element group 49: 	 $exit
      -- 
    sra_i_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 25) := "sra_i_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= sra_i_CP_1389_elements(5) & sra_i_CP_1389_elements(30) & sra_i_CP_1389_elements(33) & sra_i_CP_1389_elements(38) & sra_i_CP_1389_elements(40);
      gj_sra_i_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sra_i_CP_1389_elements(49), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_right_shift_403_data_0 : std_logic_vector(31 downto 0);
    signal LOAD_right_shift_403_wire : std_logic_vector(31 downto 0);
    signal LOAD_right_shift_403_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_right_shift_408_data_0 : std_logic_vector(31 downto 0);
    signal LOAD_right_shift_408_wire : std_logic_vector(31 downto 0);
    signal LOAD_right_shift_408_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_right_shift_423_data_0 : std_logic_vector(31 downto 0);
    signal LOAD_right_shift_423_wire : std_logic_vector(31 downto 0);
    signal LOAD_right_shift_423_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_right_shift_432_data_0 : std_logic_vector(31 downto 0);
    signal LOAD_right_shift_432_word_address_0 : std_logic_vector(0 downto 0);
    signal LSHR_u32_u32_385_wire : std_logic_vector(31 downto 0);
    signal MUX_393_wire : std_logic_vector(31 downto 0);
    signal MUX_399_wire : std_logic_vector(31 downto 0);
    signal NOT_u32_u32_410_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_425_wire : std_logic_vector(31 downto 0);
    signal STORE_right_shift_382_data_0 : std_logic_vector(31 downto 0);
    signal STORE_right_shift_382_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_right_shift_422_data_0 : std_logic_vector(31 downto 0);
    signal STORE_right_shift_422_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_right_shift_428_data_0 : std_logic_vector(31 downto 0);
    signal STORE_right_shift_428_word_address_0 : std_logic_vector(0 downto 0);
    signal SUB_u32_u32_418_wire : std_logic_vector(31 downto 0);
    signal UGT_u32_u1_396_wire : std_logic_vector(0 downto 0);
    signal ULT_u32_u1_390_wire : std_logic_vector(0 downto 0);
    signal dummy_438 : std_logic_vector(31 downto 0);
    signal konst_389_wire_constant : std_logic_vector(31 downto 0);
    signal konst_391_wire_constant : std_logic_vector(31 downto 0);
    signal konst_392_wire_constant : std_logic_vector(31 downto 0);
    signal konst_395_wire_constant : std_logic_vector(31 downto 0);
    signal konst_397_wire_constant : std_logic_vector(31 downto 0);
    signal konst_398_wire_constant : std_logic_vector(31 downto 0);
    signal konst_415_wire_constant : std_logic_vector(31 downto 0);
    signal konst_416_wire_constant : std_logic_vector(31 downto 0);
    signal konst_429_wire_constant : std_logic_vector(31 downto 0);
    signal konst_434_wire_constant : std_logic_vector(0 downto 0);
    signal konst_441_wire_constant : std_logic_vector(7 downto 0);
    signal new_420 : std_logic_vector(31 downto 0);
    signal no_of_shifts_401 : std_logic_vector(31 downto 0);
    signal output_433 : std_logic_vector(31 downto 0);
    signal sraa_406 : std_logic_vector(31 downto 0);
    signal sraaa_412 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_right_shift_403_word_address_0 <= "0";
    LOAD_right_shift_408_word_address_0 <= "0";
    LOAD_right_shift_423_word_address_0 <= "0";
    LOAD_right_shift_432_word_address_0 <= "0";
    STORE_right_shift_382_word_address_0 <= "0";
    STORE_right_shift_422_word_address_0 <= "0";
    STORE_right_shift_428_word_address_0 <= "0";
    konst_389_wire_constant <= "00000000000000000000000000100001";
    konst_391_wire_constant <= "00000000000000000000000000000001";
    konst_392_wire_constant <= "00000000000000000000000000000000";
    konst_395_wire_constant <= "00000000000000000000000000100000";
    konst_397_wire_constant <= "00000000000000000000000000000000";
    konst_398_wire_constant <= "00000000000000000000000000000000";
    konst_415_wire_constant <= "11111111111111111111111111111111";
    konst_416_wire_constant <= "00000000000000000000000000100000";
    konst_429_wire_constant <= "11111111111111111111111111111111";
    konst_434_wire_constant <= "0";
    konst_441_wire_constant <= "00000001";
    -- flow-through select operator MUX_393_inst
    MUX_393_wire <= konst_391_wire_constant when (ULT_u32_u1_390_wire(0) /=  '0') else konst_392_wire_constant;
    -- flow-through select operator MUX_399_inst
    MUX_399_wire <= konst_397_wire_constant when (UGT_u32_u1_396_wire(0) /=  '0') else konst_398_wire_constant;
    -- equivalence LOAD_right_shift_403_gather_scatter
    process(LOAD_right_shift_403_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_right_shift_403_data_0;
      ov(31 downto 0) := iv;
      LOAD_right_shift_403_wire <= ov(31 downto 0);
      --
    end process;
    -- equivalence LOAD_right_shift_408_gather_scatter
    process(LOAD_right_shift_408_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_right_shift_408_data_0;
      ov(31 downto 0) := iv;
      LOAD_right_shift_408_wire <= ov(31 downto 0);
      --
    end process;
    -- equivalence LOAD_right_shift_423_gather_scatter
    process(LOAD_right_shift_423_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_right_shift_423_data_0;
      ov(31 downto 0) := iv;
      LOAD_right_shift_423_wire <= ov(31 downto 0);
      --
    end process;
    -- equivalence LOAD_right_shift_432_gather_scatter
    process(LOAD_right_shift_432_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_right_shift_432_data_0;
      ov(31 downto 0) := iv;
      output_433 <= ov(31 downto 0);
      --
    end process;
    -- equivalence STORE_right_shift_382_gather_scatter
    process(LSHR_u32_u32_385_wire) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u32_u32_385_wire;
      ov(31 downto 0) := iv;
      STORE_right_shift_382_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence STORE_right_shift_422_gather_scatter
    process(OR_u32_u32_425_wire) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := OR_u32_u32_425_wire;
      ov(31 downto 0) := iv;
      STORE_right_shift_422_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence STORE_right_shift_428_gather_scatter
    process(konst_429_wire_constant) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := konst_429_wire_constant;
      ov(31 downto 0) := iv;
      STORE_right_shift_428_data_0 <= ov(31 downto 0);
      --
    end process;
    -- shared split operator group (0) : ADD_u8_u8_442_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pc_buffer;
      next_pc_buffer <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_442_inst_req_0;
      ADD_u8_u8_442_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_442_inst_req_1;
      ADD_u8_u8_442_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : AND_u32_u32_405_inst 
    ApIntAnd_group_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LOAD_right_shift_403_wire & no_of_shifts_401;
      sraa_406 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_405_inst_req_0;
      AND_u32_u32_405_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_405_inst_req_1;
      AND_u32_u32_405_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : AND_u32_u32_411_inst 
    ApIntAnd_group_2: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LOAD_right_shift_408_wire & NOT_u32_u32_410_wire;
      sraaa_412 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u32_u32_411_inst_req_0;
      AND_u32_u32_411_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u32_u32_411_inst_req_1;
      AND_u32_u32_411_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_2_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : LSHR_u32_u32_385_inst 
    ApIntLSHR_group_3: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= rs1_data_buffer & rs2_data_buffer;
      LSHR_u32_u32_385_wire <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_385_inst_req_0;
      LSHR_u32_u32_385_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_385_inst_req_1;
      LSHR_u32_u32_385_inst_ack_1 <= ackR_unguarded(0);
      ApIntLSHR_group_3_gI: SplitGuardInterface generic map(name => "ApIntLSHR_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- unary operator NOT_u32_u32_410_inst
    process(no_of_shifts_401) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", no_of_shifts_401, tmp_var);
      NOT_u32_u32_410_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (5) : OR_u32_u32_400_inst 
    ApIntOr_group_5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= MUX_393_wire & MUX_399_wire;
      no_of_shifts_401 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u32_u32_400_inst_req_0;
      OR_u32_u32_400_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_400_inst_req_1;
      OR_u32_u32_400_inst_ack_1 <= ackR_unguarded(0);
      ApIntOr_group_5_gI: SplitGuardInterface generic map(name => "ApIntOr_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : OR_u32_u32_425_inst 
    ApIntOr_group_6: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LOAD_right_shift_423_wire & new_420;
      OR_u32_u32_425_wire <= data_out(31 downto 0);
      guard_vector(0)  <= sraa_406(0);
      reqL_unguarded(0) <= OR_u32_u32_425_inst_req_0;
      OR_u32_u32_425_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u32_u32_425_inst_req_1;
      OR_u32_u32_425_inst_ack_1 <= ackR_unguarded(0);
      ApIntOr_group_6_gI: SplitGuardInterface generic map(name => "ApIntOr_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : SHL_u32_u32_419_inst 
    ApIntSHL_group_7: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= konst_415_wire_constant & SUB_u32_u32_418_wire;
      new_420 <= data_out(31 downto 0);
      guard_vector(0)  <= sraa_406(0);
      reqL_unguarded(0) <= SHL_u32_u32_419_inst_req_0;
      SHL_u32_u32_419_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SHL_u32_u32_419_inst_req_1;
      SHL_u32_u32_419_inst_ack_1 <= ackR_unguarded(0);
      ApIntSHL_group_7_gI: SplitGuardInterface generic map(name => "ApIntSHL_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          name => "ApIntSHL_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- binary operator SUB_u32_u32_418_inst
    process(konst_416_wire_constant, rs1_data_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_416_wire_constant, rs1_data_buffer, tmp_var);
      SUB_u32_u32_418_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_396_inst
    process(rs2_data_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(rs2_data_buffer, konst_395_wire_constant, tmp_var);
      UGT_u32_u1_396_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_390_inst
    process(rs2_data_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(rs2_data_buffer, konst_389_wire_constant, tmp_var);
      ULT_u32_u1_390_wire <= tmp_var; --
    end process;
    -- shared load operator group (0) : LOAD_right_shift_403_load_0 LOAD_right_shift_408_load_0 LOAD_right_shift_423_load_0 LOAD_right_shift_432_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => true, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      reqL_unguarded(3) <= LOAD_right_shift_403_load_0_req_0;
      reqL_unguarded(2) <= LOAD_right_shift_408_load_0_req_0;
      reqL_unguarded(1) <= LOAD_right_shift_423_load_0_req_0;
      reqL_unguarded(0) <= LOAD_right_shift_432_load_0_req_0;
      LOAD_right_shift_403_load_0_ack_0 <= ackL_unguarded(3);
      LOAD_right_shift_408_load_0_ack_0 <= ackL_unguarded(2);
      LOAD_right_shift_423_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_right_shift_432_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= LOAD_right_shift_403_load_0_req_1;
      reqR_unguarded(2) <= LOAD_right_shift_408_load_0_req_1;
      reqR_unguarded(1) <= LOAD_right_shift_423_load_0_req_1;
      reqR_unguarded(0) <= LOAD_right_shift_432_load_0_req_1;
      LOAD_right_shift_403_load_0_ack_1 <= ackR_unguarded(3);
      LOAD_right_shift_408_load_0_ack_1 <= ackR_unguarded(2);
      LOAD_right_shift_423_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_right_shift_432_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <= sraa_406(0);
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_right_shift_403_word_address_0 & LOAD_right_shift_408_word_address_0 & LOAD_right_shift_423_word_address_0 & LOAD_right_shift_432_word_address_0;
      LOAD_right_shift_403_data_0 <= data_out(127 downto 96);
      LOAD_right_shift_408_data_0 <= data_out(95 downto 64);
      LOAD_right_shift_423_data_0 <= data_out(63 downto 32);
      LOAD_right_shift_432_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(0 downto 0),
          mtag => memory_space_3_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : STORE_right_shift_382_store_0 STORE_right_shift_422_store_0 STORE_right_shift_428_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(2 downto 0);
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => true, 1 => true, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= STORE_right_shift_382_store_0_req_0;
      reqL_unguarded(1) <= STORE_right_shift_422_store_0_req_0;
      reqL_unguarded(0) <= STORE_right_shift_428_store_0_req_0;
      STORE_right_shift_382_store_0_ack_0 <= ackL_unguarded(2);
      STORE_right_shift_422_store_0_ack_0 <= ackL_unguarded(1);
      STORE_right_shift_428_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= STORE_right_shift_382_store_0_req_1;
      reqR_unguarded(1) <= STORE_right_shift_422_store_0_req_1;
      reqR_unguarded(0) <= STORE_right_shift_428_store_0_req_1;
      STORE_right_shift_382_store_0_ack_1 <= ackR_unguarded(2);
      STORE_right_shift_422_store_0_ack_1 <= ackR_unguarded(1);
      STORE_right_shift_428_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= sraaa_412(0);
      guard_vector(1)  <= sraa_406(0);
      guard_vector(2)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_right_shift_382_word_address_0 & STORE_right_shift_422_word_address_0 & STORE_right_shift_428_word_address_0;
      data_in <= STORE_right_shift_382_data_0 & STORE_right_shift_422_data_0 & STORE_right_shift_428_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 32,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(0 downto 0),
          mdata => memory_space_3_sr_data(31 downto 0),
          mtag => memory_space_3_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 3,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared call operator group (0) : call_stmt_438_call 
    accessreg_call_group_0: Block -- 
      signal data_in: std_logic_vector(40 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_438_call_req_0;
      call_stmt_438_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_438_call_req_1;
      call_stmt_438_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessreg_call_group_0_gI: SplitGuardInterface generic map(name => "accessreg_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_434_wire_constant & rd_buffer & output_433;
      dummy_438 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 41,
        owidth => 41,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessreg_call_reqs(0),
          ackR => accessreg_call_acks(0),
          dataR => accessreg_call_data(40 downto 0),
          tagR => accessreg_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessreg_return_acks(0), -- cross-over
          ackL => accessreg_return_reqs(0), -- cross-over
          dataL => accessreg_return_data(31 downto 0),
          tagL => accessreg_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end sra_i_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity srl_i is -- 
  generic (tag_length : integer); 
  port ( -- 
    rs1_data : in  std_logic_vector(31 downto 0);
    rs2_data : in  std_logic_vector(31 downto 0);
    rd : in  std_logic_vector(7 downto 0);
    pc : in  std_logic_vector(7 downto 0);
    next_pc : out  std_logic_vector(7 downto 0);
    accessreg_call_reqs : out  std_logic_vector(0 downto 0);
    accessreg_call_acks : in   std_logic_vector(0 downto 0);
    accessreg_call_data : out  std_logic_vector(40 downto 0);
    accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
    accessreg_return_reqs : out  std_logic_vector(0 downto 0);
    accessreg_return_acks : in   std_logic_vector(0 downto 0);
    accessreg_return_data : in   std_logic_vector(31 downto 0);
    accessreg_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity srl_i;
architecture srl_i_arch of srl_i is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 80)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rs1_data_buffer :  std_logic_vector(31 downto 0);
  signal rs1_data_update_enable: Boolean;
  signal rs2_data_buffer :  std_logic_vector(31 downto 0);
  signal rs2_data_update_enable: Boolean;
  signal rd_buffer :  std_logic_vector(7 downto 0);
  signal rd_update_enable: Boolean;
  signal pc_buffer :  std_logic_vector(7 downto 0);
  signal pc_update_enable: Boolean;
  -- output port buffer signals
  signal next_pc_buffer :  std_logic_vector(7 downto 0);
  signal next_pc_update_enable: Boolean;
  signal srl_i_CP_1746_start: Boolean;
  signal srl_i_CP_1746_symbol: Boolean;
  -- volatile/operator module components. 
  component accessreg is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(7 downto 0);
      write_data : in  std_logic_vector(31 downto 0);
      read_data : out  std_logic_vector(31 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal LSHR_u32_u32_454_inst_req_0 : boolean;
  signal LSHR_u32_u32_454_inst_ack_0 : boolean;
  signal LSHR_u32_u32_454_inst_req_1 : boolean;
  signal LSHR_u32_u32_454_inst_ack_1 : boolean;
  signal call_stmt_460_call_req_0 : boolean;
  signal call_stmt_460_call_ack_0 : boolean;
  signal call_stmt_460_call_req_1 : boolean;
  signal call_stmt_460_call_ack_1 : boolean;
  signal ADD_u8_u8_464_inst_req_0 : boolean;
  signal ADD_u8_u8_464_inst_ack_0 : boolean;
  signal ADD_u8_u8_464_inst_req_1 : boolean;
  signal ADD_u8_u8_464_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "srl_i_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 80) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= rs1_data;
  rs1_data_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= rs2_data;
  rs2_data_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(71 downto 64) <= rd;
  rd_buffer <= in_buffer_data_out(71 downto 64);
  in_buffer_data_in(79 downto 72) <= pc;
  pc_buffer <= in_buffer_data_out(79 downto 72);
  in_buffer_data_in(tag_length + 79 downto 80) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 79 downto 80);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  srl_i_CP_1746_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "srl_i_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= next_pc_buffer;
  next_pc <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= srl_i_CP_1746_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= srl_i_CP_1746_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= srl_i_CP_1746_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  srl_i_CP_1746: Block -- control-path 
    signal srl_i_CP_1746_elements: BooleanArray(7 downto 0);
    -- 
  begin -- 
    srl_i_CP_1746_elements(0) <= srl_i_CP_1746_start;
    srl_i_CP_1746_symbol <= srl_i_CP_1746_elements(7);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (17) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_455_to_assign_stmt_465/$entry
      -- CP-element group 0: 	 assign_stmt_455_to_assign_stmt_465/LSHR_u32_u32_454_sample_start_
      -- CP-element group 0: 	 assign_stmt_455_to_assign_stmt_465/LSHR_u32_u32_454_update_start_
      -- CP-element group 0: 	 assign_stmt_455_to_assign_stmt_465/LSHR_u32_u32_454_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_455_to_assign_stmt_465/LSHR_u32_u32_454_Sample/rr
      -- CP-element group 0: 	 assign_stmt_455_to_assign_stmt_465/LSHR_u32_u32_454_Update/$entry
      -- CP-element group 0: 	 assign_stmt_455_to_assign_stmt_465/LSHR_u32_u32_454_Update/cr
      -- CP-element group 0: 	 assign_stmt_455_to_assign_stmt_465/call_stmt_460_update_start_
      -- CP-element group 0: 	 assign_stmt_455_to_assign_stmt_465/call_stmt_460_Update/$entry
      -- CP-element group 0: 	 assign_stmt_455_to_assign_stmt_465/call_stmt_460_Update/ccr
      -- CP-element group 0: 	 assign_stmt_455_to_assign_stmt_465/ADD_u8_u8_464_sample_start_
      -- CP-element group 0: 	 assign_stmt_455_to_assign_stmt_465/ADD_u8_u8_464_update_start_
      -- CP-element group 0: 	 assign_stmt_455_to_assign_stmt_465/ADD_u8_u8_464_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_455_to_assign_stmt_465/ADD_u8_u8_464_Sample/rr
      -- CP-element group 0: 	 assign_stmt_455_to_assign_stmt_465/ADD_u8_u8_464_Update/$entry
      -- CP-element group 0: 	 assign_stmt_455_to_assign_stmt_465/ADD_u8_u8_464_Update/cr
      -- 
    ccr_1778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => srl_i_CP_1746_elements(0), ack => call_stmt_460_call_req_1); -- 
    rr_1787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => srl_i_CP_1746_elements(0), ack => ADD_u8_u8_464_inst_req_0); -- 
    cr_1792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => srl_i_CP_1746_elements(0), ack => ADD_u8_u8_464_inst_req_1); -- 
    rr_1759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => srl_i_CP_1746_elements(0), ack => LSHR_u32_u32_454_inst_req_0); -- 
    cr_1764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => srl_i_CP_1746_elements(0), ack => LSHR_u32_u32_454_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_455_to_assign_stmt_465/LSHR_u32_u32_454_sample_completed_
      -- CP-element group 1: 	 assign_stmt_455_to_assign_stmt_465/LSHR_u32_u32_454_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_455_to_assign_stmt_465/LSHR_u32_u32_454_Sample/ra
      -- 
    ra_1760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_454_inst_ack_0, ack => srl_i_CP_1746_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_455_to_assign_stmt_465/LSHR_u32_u32_454_update_completed_
      -- CP-element group 2: 	 assign_stmt_455_to_assign_stmt_465/LSHR_u32_u32_454_Update/$exit
      -- CP-element group 2: 	 assign_stmt_455_to_assign_stmt_465/LSHR_u32_u32_454_Update/ca
      -- CP-element group 2: 	 assign_stmt_455_to_assign_stmt_465/call_stmt_460_sample_start_
      -- CP-element group 2: 	 assign_stmt_455_to_assign_stmt_465/call_stmt_460_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_455_to_assign_stmt_465/call_stmt_460_Sample/crr
      -- 
    ca_1765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LSHR_u32_u32_454_inst_ack_1, ack => srl_i_CP_1746_elements(2)); -- 
    crr_1773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => srl_i_CP_1746_elements(2), ack => call_stmt_460_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_455_to_assign_stmt_465/call_stmt_460_sample_completed_
      -- CP-element group 3: 	 assign_stmt_455_to_assign_stmt_465/call_stmt_460_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_455_to_assign_stmt_465/call_stmt_460_Sample/cra
      -- 
    cra_1774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_460_call_ack_0, ack => srl_i_CP_1746_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_455_to_assign_stmt_465/call_stmt_460_update_completed_
      -- CP-element group 4: 	 assign_stmt_455_to_assign_stmt_465/call_stmt_460_Update/$exit
      -- CP-element group 4: 	 assign_stmt_455_to_assign_stmt_465/call_stmt_460_Update/cca
      -- 
    cca_1779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_460_call_ack_1, ack => srl_i_CP_1746_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_455_to_assign_stmt_465/ADD_u8_u8_464_sample_completed_
      -- CP-element group 5: 	 assign_stmt_455_to_assign_stmt_465/ADD_u8_u8_464_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_455_to_assign_stmt_465/ADD_u8_u8_464_Sample/ra
      -- 
    ra_1788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_464_inst_ack_0, ack => srl_i_CP_1746_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_455_to_assign_stmt_465/ADD_u8_u8_464_update_completed_
      -- CP-element group 6: 	 assign_stmt_455_to_assign_stmt_465/ADD_u8_u8_464_Update/$exit
      -- CP-element group 6: 	 assign_stmt_455_to_assign_stmt_465/ADD_u8_u8_464_Update/ca
      -- 
    ca_1793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_464_inst_ack_1, ack => srl_i_CP_1746_elements(6)); -- 
    -- CP-element group 7:  join  transition  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 $exit
      -- CP-element group 7: 	 assign_stmt_455_to_assign_stmt_465/$exit
      -- 
    srl_i_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "srl_i_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= srl_i_CP_1746_elements(4) & srl_i_CP_1746_elements(6);
      gj_srl_i_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => srl_i_CP_1746_elements(7), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal dummy_460 : std_logic_vector(31 downto 0);
    signal konst_456_wire_constant : std_logic_vector(0 downto 0);
    signal konst_463_wire_constant : std_logic_vector(7 downto 0);
    signal output_455 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_456_wire_constant <= "0";
    konst_463_wire_constant <= "00000001";
    -- shared split operator group (0) : ADD_u8_u8_464_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pc_buffer;
      next_pc_buffer <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_464_inst_req_0;
      ADD_u8_u8_464_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_464_inst_req_1;
      ADD_u8_u8_464_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : LSHR_u32_u32_454_inst 
    ApIntLSHR_group_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= rs1_data_buffer & rs2_data_buffer;
      output_455 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= LSHR_u32_u32_454_inst_req_0;
      LSHR_u32_u32_454_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LSHR_u32_u32_454_inst_req_1;
      LSHR_u32_u32_454_inst_ack_1 <= ackR_unguarded(0);
      ApIntLSHR_group_1_gI: SplitGuardInterface generic map(name => "ApIntLSHR_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          name => "ApIntLSHR_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared call operator group (0) : call_stmt_460_call 
    accessreg_call_group_0: Block -- 
      signal data_in: std_logic_vector(40 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_460_call_req_0;
      call_stmt_460_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_460_call_req_1;
      call_stmt_460_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessreg_call_group_0_gI: SplitGuardInterface generic map(name => "accessreg_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_456_wire_constant & rd_buffer & output_455;
      dummy_460 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 41,
        owidth => 41,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessreg_call_reqs(0),
          ackR => accessreg_call_acks(0),
          dataR => accessreg_call_data(40 downto 0),
          tagR => accessreg_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessreg_return_acks(0), -- cross-over
          ackL => accessreg_return_reqs(0), -- cross-over
          dataL => accessreg_return_data(31 downto 0),
          tagL => accessreg_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end srl_i_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity store is -- 
  generic (tag_length : integer); 
  port ( -- 
    rs1_data : in  std_logic_vector(31 downto 0);
    rs2_data : in  std_logic_vector(31 downto 0);
    pc : in  std_logic_vector(7 downto 0);
    next_pc : out  std_logic_vector(7 downto 0);
    accessMem_call_reqs : out  std_logic_vector(0 downto 0);
    accessMem_call_acks : in   std_logic_vector(0 downto 0);
    accessMem_call_data : out  std_logic_vector(40 downto 0);
    accessMem_call_tag  :  out  std_logic_vector(0 downto 0);
    accessMem_return_reqs : out  std_logic_vector(0 downto 0);
    accessMem_return_acks : in   std_logic_vector(0 downto 0);
    accessMem_return_data : in   std_logic_vector(31 downto 0);
    accessMem_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity store;
architecture store_arch of store is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 72)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rs1_data_buffer :  std_logic_vector(31 downto 0);
  signal rs1_data_update_enable: Boolean;
  signal rs2_data_buffer :  std_logic_vector(31 downto 0);
  signal rs2_data_update_enable: Boolean;
  signal pc_buffer :  std_logic_vector(7 downto 0);
  signal pc_update_enable: Boolean;
  -- output port buffer signals
  signal next_pc_buffer :  std_logic_vector(7 downto 0);
  signal next_pc_update_enable: Boolean;
  signal store_CP_1794_start: Boolean;
  signal store_CP_1794_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(7 downto 0);
      write_data : in  std_logic_vector(31 downto 0);
      read_data : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_480_call_req_1 : boolean;
  signal ADD_u8_u8_484_inst_ack_1 : boolean;
  signal ADD_u8_u8_484_inst_req_1 : boolean;
  signal call_stmt_480_call_ack_1 : boolean;
  signal ADD_u8_u8_484_inst_req_0 : boolean;
  signal call_stmt_480_call_req_0 : boolean;
  signal ADD_u8_u8_484_inst_ack_0 : boolean;
  signal call_stmt_480_call_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "store_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 72) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= rs1_data;
  rs1_data_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= rs2_data;
  rs2_data_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(71 downto 64) <= pc;
  pc_buffer <= in_buffer_data_out(71 downto 64);
  in_buffer_data_in(tag_length + 71 downto 72) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 71 downto 72);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  store_CP_1794_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "store_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= next_pc_buffer;
  next_pc <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= store_CP_1794_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= store_CP_1794_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= store_CP_1794_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  store_CP_1794: Block -- control-path 
    signal store_CP_1794_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    store_CP_1794_elements(0) <= store_CP_1794_start;
    store_CP_1794_symbol <= store_CP_1794_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 assign_stmt_475_to_assign_stmt_485/call_stmt_480_Update/ccr
      -- CP-element group 0: 	 assign_stmt_475_to_assign_stmt_485/ADD_u8_u8_484_Update/$entry
      -- CP-element group 0: 	 assign_stmt_475_to_assign_stmt_485/call_stmt_480_Update/$entry
      -- CP-element group 0: 	 assign_stmt_475_to_assign_stmt_485/ADD_u8_u8_484_sample_start_
      -- CP-element group 0: 	 assign_stmt_475_to_assign_stmt_485/ADD_u8_u8_484_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_475_to_assign_stmt_485/$entry
      -- CP-element group 0: 	 assign_stmt_475_to_assign_stmt_485/ADD_u8_u8_484_Update/cr
      -- CP-element group 0: 	 assign_stmt_475_to_assign_stmt_485/ADD_u8_u8_484_update_start_
      -- CP-element group 0: 	 assign_stmt_475_to_assign_stmt_485/call_stmt_480_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_475_to_assign_stmt_485/ADD_u8_u8_484_Sample/rr
      -- CP-element group 0: 	 assign_stmt_475_to_assign_stmt_485/call_stmt_480_Sample/crr
      -- CP-element group 0: 	 assign_stmt_475_to_assign_stmt_485/call_stmt_480_sample_start_
      -- CP-element group 0: 	 assign_stmt_475_to_assign_stmt_485/call_stmt_480_update_start_
      -- CP-element group 0: 	 $entry
      -- 
    crr_1807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => store_CP_1794_elements(0), ack => call_stmt_480_call_req_0); -- 
    ccr_1812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => store_CP_1794_elements(0), ack => call_stmt_480_call_req_1); -- 
    rr_1821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => store_CP_1794_elements(0), ack => ADD_u8_u8_484_inst_req_0); -- 
    cr_1826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => store_CP_1794_elements(0), ack => ADD_u8_u8_484_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_475_to_assign_stmt_485/call_stmt_480_Sample/cra
      -- CP-element group 1: 	 assign_stmt_475_to_assign_stmt_485/call_stmt_480_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_475_to_assign_stmt_485/call_stmt_480_sample_completed_
      -- 
    cra_1808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_480_call_ack_0, ack => store_CP_1794_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_475_to_assign_stmt_485/call_stmt_480_Update/cca
      -- CP-element group 2: 	 assign_stmt_475_to_assign_stmt_485/call_stmt_480_Update/$exit
      -- CP-element group 2: 	 assign_stmt_475_to_assign_stmt_485/call_stmt_480_update_completed_
      -- 
    cca_1813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_480_call_ack_1, ack => store_CP_1794_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_475_to_assign_stmt_485/ADD_u8_u8_484_Sample/ra
      -- CP-element group 3: 	 assign_stmt_475_to_assign_stmt_485/ADD_u8_u8_484_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_475_to_assign_stmt_485/ADD_u8_u8_484_sample_completed_
      -- 
    ra_1822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_484_inst_ack_0, ack => store_CP_1794_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_475_to_assign_stmt_485/ADD_u8_u8_484_update_completed_
      -- CP-element group 4: 	 assign_stmt_475_to_assign_stmt_485/ADD_u8_u8_484_Update/ca
      -- CP-element group 4: 	 assign_stmt_475_to_assign_stmt_485/ADD_u8_u8_484_Update/$exit
      -- 
    ca_1827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_484_inst_ack_1, ack => store_CP_1794_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_475_to_assign_stmt_485/$exit
      -- CP-element group 5: 	 $exit
      -- 
    store_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "store_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= store_CP_1794_elements(2) & store_CP_1794_elements(4);
      gj_store_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => store_CP_1794_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal addr_475 : std_logic_vector(7 downto 0);
    signal dummy1_480 : std_logic_vector(31 downto 0);
    signal konst_476_wire_constant : std_logic_vector(0 downto 0);
    signal konst_483_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_476_wire_constant <= "0";
    konst_483_wire_constant <= "00000001";
    -- flow-through slice operator slice_474_inst
    addr_475 <= rs1_data_buffer(7 downto 0);
    -- shared split operator group (0) : ADD_u8_u8_484_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pc_buffer;
      next_pc_buffer <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_484_inst_req_0;
      ADD_u8_u8_484_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_484_inst_req_1;
      ADD_u8_u8_484_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared call operator group (0) : call_stmt_480_call 
    accessMem_call_group_0: Block -- 
      signal data_in: std_logic_vector(40 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_480_call_req_0;
      call_stmt_480_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_480_call_req_1;
      call_stmt_480_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMem_call_group_0_gI: SplitGuardInterface generic map(name => "accessMem_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_476_wire_constant & addr_475 & rs2_data_buffer;
      dummy1_480 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 41,
        owidth => 41,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMem_call_reqs(0),
          ackR => accessMem_call_acks(0),
          dataR => accessMem_call_data(40 downto 0),
          tagR => accessMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMem_return_acks(0), -- cross-over
          ackL => accessMem_return_reqs(0), -- cross-over
          dataL => accessMem_return_data(31 downto 0),
          tagL => accessMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end store_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sub is -- 
  generic (tag_length : integer); 
  port ( -- 
    rs1_data : in  std_logic_vector(31 downto 0);
    rs2_data : in  std_logic_vector(31 downto 0);
    rd : in  std_logic_vector(7 downto 0);
    pc : in  std_logic_vector(7 downto 0);
    next_pc : out  std_logic_vector(7 downto 0);
    accessreg_call_reqs : out  std_logic_vector(0 downto 0);
    accessreg_call_acks : in   std_logic_vector(0 downto 0);
    accessreg_call_data : out  std_logic_vector(40 downto 0);
    accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
    accessreg_return_reqs : out  std_logic_vector(0 downto 0);
    accessreg_return_acks : in   std_logic_vector(0 downto 0);
    accessreg_return_data : in   std_logic_vector(31 downto 0);
    accessreg_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sub;
architecture sub_arch of sub is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 80)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rs1_data_buffer :  std_logic_vector(31 downto 0);
  signal rs1_data_update_enable: Boolean;
  signal rs2_data_buffer :  std_logic_vector(31 downto 0);
  signal rs2_data_update_enable: Boolean;
  signal rd_buffer :  std_logic_vector(7 downto 0);
  signal rd_update_enable: Boolean;
  signal pc_buffer :  std_logic_vector(7 downto 0);
  signal pc_update_enable: Boolean;
  -- output port buffer signals
  signal next_pc_buffer :  std_logic_vector(7 downto 0);
  signal next_pc_update_enable: Boolean;
  signal sub_CP_1828_start: Boolean;
  signal sub_CP_1828_symbol: Boolean;
  -- volatile/operator module components. 
  component accessreg is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(7 downto 0);
      write_data : in  std_logic_vector(31 downto 0);
      read_data : out  std_logic_vector(31 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal ADD_u8_u8_506_inst_req_1 : boolean;
  signal call_stmt_502_call_ack_1 : boolean;
  signal call_stmt_502_call_req_1 : boolean;
  signal ADD_u8_u8_506_inst_ack_1 : boolean;
  signal call_stmt_502_call_ack_0 : boolean;
  signal call_stmt_502_call_req_0 : boolean;
  signal ADD_u8_u8_506_inst_ack_0 : boolean;
  signal SUB_u32_u32_496_inst_ack_1 : boolean;
  signal SUB_u32_u32_496_inst_req_1 : boolean;
  signal ADD_u8_u8_506_inst_req_0 : boolean;
  signal SUB_u32_u32_496_inst_ack_0 : boolean;
  signal SUB_u32_u32_496_inst_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sub_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 80) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= rs1_data;
  rs1_data_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= rs2_data;
  rs2_data_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(71 downto 64) <= rd;
  rd_buffer <= in_buffer_data_out(71 downto 64);
  in_buffer_data_in(79 downto 72) <= pc;
  pc_buffer <= in_buffer_data_out(79 downto 72);
  in_buffer_data_in(tag_length + 79 downto 80) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 79 downto 80);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sub_CP_1828_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sub_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= next_pc_buffer;
  next_pc <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sub_CP_1828_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sub_CP_1828_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sub_CP_1828_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sub_CP_1828: Block -- control-path 
    signal sub_CP_1828_elements: BooleanArray(7 downto 0);
    -- 
  begin -- 
    sub_CP_1828_elements(0) <= sub_CP_1828_start;
    sub_CP_1828_symbol <= sub_CP_1828_elements(7);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (17) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_497_to_assign_stmt_507/ADD_u8_u8_506_Update/cr
      -- CP-element group 0: 	 assign_stmt_497_to_assign_stmt_507/$entry
      -- CP-element group 0: 	 assign_stmt_497_to_assign_stmt_507/call_stmt_502_Update/ccr
      -- CP-element group 0: 	 assign_stmt_497_to_assign_stmt_507/call_stmt_502_Update/$entry
      -- CP-element group 0: 	 assign_stmt_497_to_assign_stmt_507/call_stmt_502_update_start_
      -- CP-element group 0: 	 assign_stmt_497_to_assign_stmt_507/ADD_u8_u8_506_Update/$entry
      -- CP-element group 0: 	 assign_stmt_497_to_assign_stmt_507/SUB_u32_u32_496_sample_start_
      -- CP-element group 0: 	 assign_stmt_497_to_assign_stmt_507/ADD_u8_u8_506_sample_start_
      -- CP-element group 0: 	 assign_stmt_497_to_assign_stmt_507/ADD_u8_u8_506_update_start_
      -- CP-element group 0: 	 assign_stmt_497_to_assign_stmt_507/SUB_u32_u32_496_update_start_
      -- CP-element group 0: 	 assign_stmt_497_to_assign_stmt_507/SUB_u32_u32_496_Update/cr
      -- CP-element group 0: 	 assign_stmt_497_to_assign_stmt_507/ADD_u8_u8_506_Sample/rr
      -- CP-element group 0: 	 assign_stmt_497_to_assign_stmt_507/SUB_u32_u32_496_Update/$entry
      -- CP-element group 0: 	 assign_stmt_497_to_assign_stmt_507/SUB_u32_u32_496_Sample/rr
      -- CP-element group 0: 	 assign_stmt_497_to_assign_stmt_507/SUB_u32_u32_496_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_497_to_assign_stmt_507/ADD_u8_u8_506_Sample/$entry
      -- 
    cr_1846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sub_CP_1828_elements(0), ack => SUB_u32_u32_496_inst_req_1); -- 
    rr_1869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sub_CP_1828_elements(0), ack => ADD_u8_u8_506_inst_req_0); -- 
    cr_1874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sub_CP_1828_elements(0), ack => ADD_u8_u8_506_inst_req_1); -- 
    ccr_1860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sub_CP_1828_elements(0), ack => call_stmt_502_call_req_1); -- 
    rr_1841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sub_CP_1828_elements(0), ack => SUB_u32_u32_496_inst_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_497_to_assign_stmt_507/SUB_u32_u32_496_sample_completed_
      -- CP-element group 1: 	 assign_stmt_497_to_assign_stmt_507/SUB_u32_u32_496_Sample/ra
      -- CP-element group 1: 	 assign_stmt_497_to_assign_stmt_507/SUB_u32_u32_496_Sample/$exit
      -- 
    ra_1842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_496_inst_ack_0, ack => sub_CP_1828_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_497_to_assign_stmt_507/call_stmt_502_Sample/crr
      -- CP-element group 2: 	 assign_stmt_497_to_assign_stmt_507/call_stmt_502_sample_start_
      -- CP-element group 2: 	 assign_stmt_497_to_assign_stmt_507/SUB_u32_u32_496_Update/ca
      -- CP-element group 2: 	 assign_stmt_497_to_assign_stmt_507/call_stmt_502_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_497_to_assign_stmt_507/SUB_u32_u32_496_Update/$exit
      -- CP-element group 2: 	 assign_stmt_497_to_assign_stmt_507/SUB_u32_u32_496_update_completed_
      -- 
    ca_1847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_496_inst_ack_1, ack => sub_CP_1828_elements(2)); -- 
    crr_1855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sub_CP_1828_elements(2), ack => call_stmt_502_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_497_to_assign_stmt_507/call_stmt_502_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_497_to_assign_stmt_507/call_stmt_502_Sample/cra
      -- CP-element group 3: 	 assign_stmt_497_to_assign_stmt_507/call_stmt_502_sample_completed_
      -- 
    cra_1856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_502_call_ack_0, ack => sub_CP_1828_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_497_to_assign_stmt_507/call_stmt_502_Update/cca
      -- CP-element group 4: 	 assign_stmt_497_to_assign_stmt_507/call_stmt_502_Update/$exit
      -- CP-element group 4: 	 assign_stmt_497_to_assign_stmt_507/call_stmt_502_update_completed_
      -- 
    cca_1861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_502_call_ack_1, ack => sub_CP_1828_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_497_to_assign_stmt_507/ADD_u8_u8_506_Sample/ra
      -- CP-element group 5: 	 assign_stmt_497_to_assign_stmt_507/ADD_u8_u8_506_sample_completed_
      -- CP-element group 5: 	 assign_stmt_497_to_assign_stmt_507/ADD_u8_u8_506_Sample/$exit
      -- 
    ra_1870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_506_inst_ack_0, ack => sub_CP_1828_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_497_to_assign_stmt_507/ADD_u8_u8_506_Update/ca
      -- CP-element group 6: 	 assign_stmt_497_to_assign_stmt_507/ADD_u8_u8_506_Update/$exit
      -- CP-element group 6: 	 assign_stmt_497_to_assign_stmt_507/ADD_u8_u8_506_update_completed_
      -- 
    ca_1875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_506_inst_ack_1, ack => sub_CP_1828_elements(6)); -- 
    -- CP-element group 7:  join  transition  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 $exit
      -- CP-element group 7: 	 assign_stmt_497_to_assign_stmt_507/$exit
      -- 
    sub_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 22) := "sub_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sub_CP_1828_elements(4) & sub_CP_1828_elements(6);
      gj_sub_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sub_CP_1828_elements(7), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal dummy_502 : std_logic_vector(31 downto 0);
    signal konst_498_wire_constant : std_logic_vector(0 downto 0);
    signal konst_505_wire_constant : std_logic_vector(7 downto 0);
    signal output_497 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_498_wire_constant <= "0";
    konst_505_wire_constant <= "00000001";
    -- shared split operator group (0) : ADD_u8_u8_506_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pc_buffer;
      next_pc_buffer <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_506_inst_req_0;
      ADD_u8_u8_506_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_506_inst_req_1;
      ADD_u8_u8_506_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : SUB_u32_u32_496_inst 
    ApIntSub_group_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= rs1_data_buffer & rs2_data_buffer;
      output_497 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_496_inst_req_0;
      SUB_u32_u32_496_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_496_inst_req_1;
      SUB_u32_u32_496_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_1_gI: SplitGuardInterface generic map(name => "ApIntSub_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared call operator group (0) : call_stmt_502_call 
    accessreg_call_group_0: Block -- 
      signal data_in: std_logic_vector(40 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_502_call_req_0;
      call_stmt_502_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_502_call_req_1;
      call_stmt_502_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessreg_call_group_0_gI: SplitGuardInterface generic map(name => "accessreg_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_498_wire_constant & rd_buffer & output_497;
      dummy_502 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 41,
        owidth => 41,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessreg_call_reqs(0),
          ackR => accessreg_call_acks(0),
          dataR => accessreg_call_data(40 downto 0),
          tagR => accessreg_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessreg_return_acks(0), -- cross-over
          ackL => accessreg_return_reqs(0), -- cross-over
          dataL => accessreg_return_data(31 downto 0),
          tagL => accessreg_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end sub_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity try is -- 
  generic (tag_length : integer); 
  port ( -- 
    pc : in  std_logic_vector(7 downto 0);
    inst : in  std_logic_vector(31 downto 0);
    next_pc : out  std_logic_vector(7 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    cmp_call_reqs : out  std_logic_vector(0 downto 0);
    cmp_call_acks : in   std_logic_vector(0 downto 0);
    cmp_call_data : out  std_logic_vector(79 downto 0);
    cmp_call_tag  :  out  std_logic_vector(0 downto 0);
    cmp_return_reqs : out  std_logic_vector(0 downto 0);
    cmp_return_acks : in   std_logic_vector(0 downto 0);
    cmp_return_data : in   std_logic_vector(7 downto 0);
    cmp_return_tag :  in   std_logic_vector(0 downto 0);
    sub_call_reqs : out  std_logic_vector(0 downto 0);
    sub_call_acks : in   std_logic_vector(0 downto 0);
    sub_call_data : out  std_logic_vector(79 downto 0);
    sub_call_tag  :  out  std_logic_vector(0 downto 0);
    sub_return_reqs : out  std_logic_vector(0 downto 0);
    sub_return_acks : in   std_logic_vector(0 downto 0);
    sub_return_data : in   std_logic_vector(7 downto 0);
    sub_return_tag :  in   std_logic_vector(0 downto 0);
    accessreg_call_reqs : out  std_logic_vector(0 downto 0);
    accessreg_call_acks : in   std_logic_vector(0 downto 0);
    accessreg_call_data : out  std_logic_vector(40 downto 0);
    accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
    accessreg_return_reqs : out  std_logic_vector(0 downto 0);
    accessreg_return_acks : in   std_logic_vector(0 downto 0);
    accessreg_return_data : in   std_logic_vector(31 downto 0);
    accessreg_return_tag :  in   std_logic_vector(1 downto 0);
    bn_call_reqs : out  std_logic_vector(0 downto 0);
    bn_call_acks : in   std_logic_vector(0 downto 0);
    bn_call_data : out  std_logic_vector(79 downto 0);
    bn_call_tag  :  out  std_logic_vector(0 downto 0);
    bn_return_reqs : out  std_logic_vector(0 downto 0);
    bn_return_acks : in   std_logic_vector(0 downto 0);
    bn_return_data : in   std_logic_vector(7 downto 0);
    bn_return_tag :  in   std_logic_vector(0 downto 0);
    halt_call_reqs : out  std_logic_vector(0 downto 0);
    halt_call_acks : in   std_logic_vector(0 downto 0);
    halt_call_data : out  std_logic_vector(7 downto 0);
    halt_call_tag  :  out  std_logic_vector(0 downto 0);
    halt_return_reqs : out  std_logic_vector(0 downto 0);
    halt_return_acks : in   std_logic_vector(0 downto 0);
    halt_return_data : in   std_logic_vector(7 downto 0);
    halt_return_tag :  in   std_logic_vector(0 downto 0);
    add_call_reqs : out  std_logic_vector(0 downto 0);
    add_call_acks : in   std_logic_vector(0 downto 0);
    add_call_data : out  std_logic_vector(79 downto 0);
    add_call_tag  :  out  std_logic_vector(0 downto 0);
    add_return_reqs : out  std_logic_vector(0 downto 0);
    add_return_acks : in   std_logic_vector(0 downto 0);
    add_return_data : in   std_logic_vector(7 downto 0);
    add_return_tag :  in   std_logic_vector(0 downto 0);
    sll_i_call_reqs : out  std_logic_vector(0 downto 0);
    sll_i_call_acks : in   std_logic_vector(0 downto 0);
    sll_i_call_data : out  std_logic_vector(79 downto 0);
    sll_i_call_tag  :  out  std_logic_vector(0 downto 0);
    sll_i_return_reqs : out  std_logic_vector(0 downto 0);
    sll_i_return_acks : in   std_logic_vector(0 downto 0);
    sll_i_return_data : in   std_logic_vector(7 downto 0);
    sll_i_return_tag :  in   std_logic_vector(0 downto 0);
    and_i_call_reqs : out  std_logic_vector(0 downto 0);
    and_i_call_acks : in   std_logic_vector(0 downto 0);
    and_i_call_data : out  std_logic_vector(79 downto 0);
    and_i_call_tag  :  out  std_logic_vector(0 downto 0);
    and_i_return_reqs : out  std_logic_vector(0 downto 0);
    and_i_return_acks : in   std_logic_vector(0 downto 0);
    and_i_return_data : in   std_logic_vector(7 downto 0);
    and_i_return_tag :  in   std_logic_vector(0 downto 0);
    call_call_reqs : out  std_logic_vector(0 downto 0);
    call_call_acks : in   std_logic_vector(0 downto 0);
    call_call_data : out  std_logic_vector(79 downto 0);
    call_call_tag  :  out  std_logic_vector(0 downto 0);
    call_return_reqs : out  std_logic_vector(0 downto 0);
    call_return_acks : in   std_logic_vector(0 downto 0);
    call_return_data : in   std_logic_vector(7 downto 0);
    call_return_tag :  in   std_logic_vector(0 downto 0);
    bz_call_reqs : out  std_logic_vector(0 downto 0);
    bz_call_acks : in   std_logic_vector(0 downto 0);
    bz_call_data : out  std_logic_vector(79 downto 0);
    bz_call_tag  :  out  std_logic_vector(0 downto 0);
    bz_return_reqs : out  std_logic_vector(0 downto 0);
    bz_return_acks : in   std_logic_vector(0 downto 0);
    bz_return_data : in   std_logic_vector(7 downto 0);
    bz_return_tag :  in   std_logic_vector(0 downto 0);
    xnor_i_call_reqs : out  std_logic_vector(0 downto 0);
    xnor_i_call_acks : in   std_logic_vector(0 downto 0);
    xnor_i_call_data : out  std_logic_vector(79 downto 0);
    xnor_i_call_tag  :  out  std_logic_vector(0 downto 0);
    xnor_i_return_reqs : out  std_logic_vector(0 downto 0);
    xnor_i_return_acks : in   std_logic_vector(0 downto 0);
    xnor_i_return_data : in   std_logic_vector(7 downto 0);
    xnor_i_return_tag :  in   std_logic_vector(0 downto 0);
    sra_i_call_reqs : out  std_logic_vector(0 downto 0);
    sra_i_call_acks : in   std_logic_vector(0 downto 0);
    sra_i_call_data : out  std_logic_vector(79 downto 0);
    sra_i_call_tag  :  out  std_logic_vector(0 downto 0);
    sra_i_return_reqs : out  std_logic_vector(0 downto 0);
    sra_i_return_acks : in   std_logic_vector(0 downto 0);
    sra_i_return_data : in   std_logic_vector(7 downto 0);
    sra_i_return_tag :  in   std_logic_vector(0 downto 0);
    sbir_call_reqs : out  std_logic_vector(0 downto 0);
    sbir_call_acks : in   std_logic_vector(0 downto 0);
    sbir_call_data : out  std_logic_vector(23 downto 0);
    sbir_call_tag  :  out  std_logic_vector(0 downto 0);
    sbir_return_reqs : out  std_logic_vector(0 downto 0);
    sbir_return_acks : in   std_logic_vector(0 downto 0);
    sbir_return_data : in   std_logic_vector(7 downto 0);
    sbir_return_tag :  in   std_logic_vector(0 downto 0);
    or_i_call_reqs : out  std_logic_vector(0 downto 0);
    or_i_call_acks : in   std_logic_vector(0 downto 0);
    or_i_call_data : out  std_logic_vector(79 downto 0);
    or_i_call_tag  :  out  std_logic_vector(0 downto 0);
    or_i_return_reqs : out  std_logic_vector(0 downto 0);
    or_i_return_acks : in   std_logic_vector(0 downto 0);
    or_i_return_data : in   std_logic_vector(7 downto 0);
    or_i_return_tag :  in   std_logic_vector(0 downto 0);
    load_call_reqs : out  std_logic_vector(0 downto 0);
    load_call_acks : in   std_logic_vector(0 downto 0);
    load_call_data : out  std_logic_vector(47 downto 0);
    load_call_tag  :  out  std_logic_vector(0 downto 0);
    load_return_reqs : out  std_logic_vector(0 downto 0);
    load_return_acks : in   std_logic_vector(0 downto 0);
    load_return_data : in   std_logic_vector(7 downto 0);
    load_return_tag :  in   std_logic_vector(0 downto 0);
    jmp_call_reqs : out  std_logic_vector(0 downto 0);
    jmp_call_acks : in   std_logic_vector(0 downto 0);
    jmp_call_data : out  std_logic_vector(39 downto 0);
    jmp_call_tag  :  out  std_logic_vector(0 downto 0);
    jmp_return_reqs : out  std_logic_vector(0 downto 0);
    jmp_return_acks : in   std_logic_vector(0 downto 0);
    jmp_return_data : in   std_logic_vector(7 downto 0);
    jmp_return_tag :  in   std_logic_vector(0 downto 0);
    store_call_reqs : out  std_logic_vector(0 downto 0);
    store_call_acks : in   std_logic_vector(0 downto 0);
    store_call_data : out  std_logic_vector(71 downto 0);
    store_call_tag  :  out  std_logic_vector(0 downto 0);
    store_return_reqs : out  std_logic_vector(0 downto 0);
    store_return_acks : in   std_logic_vector(0 downto 0);
    store_return_data : in   std_logic_vector(7 downto 0);
    store_return_tag :  in   std_logic_vector(0 downto 0);
    srl_i_call_reqs : out  std_logic_vector(0 downto 0);
    srl_i_call_acks : in   std_logic_vector(0 downto 0);
    srl_i_call_data : out  std_logic_vector(79 downto 0);
    srl_i_call_tag  :  out  std_logic_vector(0 downto 0);
    srl_i_return_reqs : out  std_logic_vector(0 downto 0);
    srl_i_return_acks : in   std_logic_vector(0 downto 0);
    srl_i_return_data : in   std_logic_vector(7 downto 0);
    srl_i_return_tag :  in   std_logic_vector(0 downto 0);
    xor_i_call_reqs : out  std_logic_vector(0 downto 0);
    xor_i_call_acks : in   std_logic_vector(0 downto 0);
    xor_i_call_data : out  std_logic_vector(79 downto 0);
    xor_i_call_tag  :  out  std_logic_vector(0 downto 0);
    xor_i_return_reqs : out  std_logic_vector(0 downto 0);
    xor_i_return_acks : in   std_logic_vector(0 downto 0);
    xor_i_return_data : in   std_logic_vector(7 downto 0);
    xor_i_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity try;
architecture try_arch of try is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 40)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal pc_buffer :  std_logic_vector(7 downto 0);
  signal pc_update_enable: Boolean;
  signal inst_buffer :  std_logic_vector(31 downto 0);
  signal inst_update_enable: Boolean;
  -- output port buffer signals
  signal next_pc_buffer :  std_logic_vector(7 downto 0);
  signal next_pc_update_enable: Boolean;
  signal try_CP_1972_start: Boolean;
  signal try_CP_1972_symbol: Boolean;
  -- volatile/operator module components. 
  component cmp is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sub is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component accessreg is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(7 downto 0);
      write_data : in  std_logic_vector(31 downto 0);
      read_data : out  std_logic_vector(31 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component bn is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component halt is -- 
    generic (tag_length : integer); 
    port ( -- 
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component add is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sll_i is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component and_i is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component call is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component bz is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component xnor_i is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sra_i is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(2 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sbir is -- 
    generic (tag_length : integer); 
    port ( -- 
      imm : in  std_logic_vector(7 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component or_i is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component load is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessMem_call_acks : in   std_logic_vector(0 downto 0);
      accessMem_call_data : out  std_logic_vector(40 downto 0);
      accessMem_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessMem_return_acks : in   std_logic_vector(0 downto 0);
      accessMem_return_data : in   std_logic_vector(31 downto 0);
      accessMem_return_tag :  in   std_logic_vector(0 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component jmp is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component store is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessMem_call_acks : in   std_logic_vector(0 downto 0);
      accessMem_call_data : out  std_logic_vector(40 downto 0);
      accessMem_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessMem_return_acks : in   std_logic_vector(0 downto 0);
      accessMem_return_data : in   std_logic_vector(31 downto 0);
      accessMem_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component srl_i is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component xor_i is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal LOAD_next_pc1_795_load_0_req_1 : boolean;
  signal LOAD_next_pc1_795_load_0_req_0 : boolean;
  signal LOAD_next_pc1_795_load_0_ack_1 : boolean;
  signal LOAD_next_pc1_795_load_0_ack_0 : boolean;
  signal call_stmt_667_call_req_0 : boolean;
  signal call_stmt_667_call_ack_0 : boolean;
  signal call_stmt_667_call_req_1 : boolean;
  signal call_stmt_667_call_ack_1 : boolean;
  signal call_stmt_672_call_req_0 : boolean;
  signal call_stmt_672_call_ack_0 : boolean;
  signal call_stmt_672_call_req_1 : boolean;
  signal call_stmt_672_call_ack_1 : boolean;
  signal call_stmt_676_call_req_0 : boolean;
  signal call_stmt_676_call_ack_0 : boolean;
  signal call_stmt_676_call_req_1 : boolean;
  signal call_stmt_676_call_ack_1 : boolean;
  signal STORE_next_pc1_675_store_0_req_0 : boolean;
  signal STORE_next_pc1_675_store_0_ack_0 : boolean;
  signal STORE_next_pc1_675_store_0_req_1 : boolean;
  signal STORE_next_pc1_675_store_0_ack_1 : boolean;
  signal call_stmt_682_call_req_0 : boolean;
  signal call_stmt_682_call_ack_0 : boolean;
  signal call_stmt_682_call_req_1 : boolean;
  signal call_stmt_682_call_ack_1 : boolean;
  signal call_stmt_688_call_req_0 : boolean;
  signal call_stmt_688_call_ack_0 : boolean;
  signal call_stmt_688_call_req_1 : boolean;
  signal call_stmt_688_call_ack_1 : boolean;
  signal call_stmt_694_call_req_0 : boolean;
  signal call_stmt_694_call_ack_0 : boolean;
  signal call_stmt_694_call_req_1 : boolean;
  signal call_stmt_694_call_ack_1 : boolean;
  signal call_stmt_701_call_req_0 : boolean;
  signal call_stmt_701_call_ack_0 : boolean;
  signal call_stmt_701_call_req_1 : boolean;
  signal call_stmt_701_call_ack_1 : boolean;
  signal call_stmt_708_call_req_0 : boolean;
  signal call_stmt_708_call_ack_0 : boolean;
  signal call_stmt_708_call_req_1 : boolean;
  signal call_stmt_708_call_ack_1 : boolean;
  signal call_stmt_715_call_req_0 : boolean;
  signal call_stmt_715_call_ack_0 : boolean;
  signal call_stmt_715_call_req_1 : boolean;
  signal call_stmt_715_call_ack_1 : boolean;
  signal call_stmt_722_call_req_0 : boolean;
  signal call_stmt_722_call_ack_0 : boolean;
  signal call_stmt_722_call_req_1 : boolean;
  signal call_stmt_722_call_ack_1 : boolean;
  signal call_stmt_729_call_req_0 : boolean;
  signal call_stmt_729_call_ack_0 : boolean;
  signal call_stmt_729_call_req_1 : boolean;
  signal call_stmt_729_call_ack_1 : boolean;
  signal call_stmt_736_call_req_0 : boolean;
  signal call_stmt_736_call_ack_0 : boolean;
  signal call_stmt_736_call_req_1 : boolean;
  signal call_stmt_736_call_ack_1 : boolean;
  signal call_stmt_743_call_req_0 : boolean;
  signal call_stmt_743_call_ack_0 : boolean;
  signal call_stmt_743_call_req_1 : boolean;
  signal call_stmt_743_call_ack_1 : boolean;
  signal call_stmt_750_call_req_0 : boolean;
  signal call_stmt_750_call_ack_0 : boolean;
  signal call_stmt_750_call_req_1 : boolean;
  signal call_stmt_750_call_ack_1 : boolean;
  signal call_stmt_757_call_req_0 : boolean;
  signal call_stmt_757_call_ack_0 : boolean;
  signal MUX_883_inst_ack_1 : boolean;
  signal call_stmt_757_call_req_1 : boolean;
  signal call_stmt_757_call_ack_1 : boolean;
  signal call_stmt_764_call_req_0 : boolean;
  signal call_stmt_764_call_ack_0 : boolean;
  signal MUX_883_inst_req_1 : boolean;
  signal call_stmt_764_call_req_1 : boolean;
  signal call_stmt_764_call_ack_1 : boolean;
  signal call_stmt_771_call_req_0 : boolean;
  signal call_stmt_771_call_ack_0 : boolean;
  signal call_stmt_771_call_req_1 : boolean;
  signal call_stmt_771_call_ack_1 : boolean;
  signal MUX_883_inst_ack_0 : boolean;
  signal call_stmt_778_call_req_0 : boolean;
  signal call_stmt_778_call_ack_0 : boolean;
  signal MUX_883_inst_req_0 : boolean;
  signal call_stmt_778_call_req_1 : boolean;
  signal call_stmt_778_call_ack_1 : boolean;
  signal call_stmt_783_call_req_0 : boolean;
  signal call_stmt_783_call_ack_0 : boolean;
  signal call_stmt_783_call_req_1 : boolean;
  signal call_stmt_783_call_ack_1 : boolean;
  signal call_stmt_790_call_req_0 : boolean;
  signal call_stmt_790_call_ack_0 : boolean;
  signal call_stmt_790_call_req_1 : boolean;
  signal call_stmt_790_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "try_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 40) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= pc;
  pc_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(39 downto 8) <= inst;
  inst_buffer <= in_buffer_data_out(39 downto 8);
  in_buffer_data_in(tag_length + 39 downto 40) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 39 downto 40);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  try_CP_1972_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "try_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= next_pc_buffer;
  next_pc <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= try_CP_1972_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= try_CP_1972_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= try_CP_1972_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  try_CP_1972: Block -- control-path 
    signal try_CP_1972_elements: BooleanArray(83 downto 0);
    -- 
  begin -- 
    try_CP_1972_elements(0) <= try_CP_1972_start;
    try_CP_1972_symbol <= try_CP_1972_elements(83);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	50 
    -- CP-element group 0: 	64 
    -- CP-element group 0: 	47 
    -- CP-element group 0: 	53 
    -- CP-element group 0: 	58 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	55 
    -- CP-element group 0: 	62 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	11 
    -- CP-element group 0: 	14 
    -- CP-element group 0: 	17 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	26 
    -- CP-element group 0: 	29 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	35 
    -- CP-element group 0: 	38 
    -- CP-element group 0: 	41 
    -- CP-element group 0: 	44 
    -- CP-element group 0:  members (85) 
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_Update/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/MUX_883_update_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_update_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_667_sample_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_667_update_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_667_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_667_Sample/crr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_667_Update/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_667_Update/ccr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_672_update_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_672_Update/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_672_Update/ccr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_676_sample_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_676_update_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_676_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_676_Sample/crr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_676_Update/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_676_Update/ccr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_update_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_Update/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_682_update_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_682_Update/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_682_Update/ccr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_688_update_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_688_Update/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_688_Update/ccr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_694_update_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_694_Update/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_694_Update/ccr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_701_update_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_701_Update/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_701_Update/ccr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_708_update_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_708_Update/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_708_Update/ccr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_715_update_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_715_Update/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_715_Update/ccr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_722_update_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_722_Update/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_722_Update/ccr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_729_update_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_729_Update/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_729_Update/ccr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_736_update_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_736_Update/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_736_Update/ccr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_743_update_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_743_Update/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_743_Update/ccr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_750_update_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_750_Update/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_750_Update/ccr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_757_update_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_757_Update/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_757_Update/ccr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_764_update_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_764_Update/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/MUX_883_complete/req
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_764_Update/ccr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_771_update_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_771_Update/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/MUX_883_complete/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_771_Update/ccr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_778_update_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_778_Update/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_778_Update/ccr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_783_update_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_783_Update/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_783_Update/ccr
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_790_update_start_
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_790_Update/$entry
      -- CP-element group 0: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_790_Update/ccr
      -- 
    ccr_1990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => call_stmt_667_call_req_1); -- 
    ccr_2004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => call_stmt_672_call_req_1); -- 
    crr_2013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => call_stmt_676_call_req_0); -- 
    ccr_2018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => call_stmt_676_call_req_1); -- 
    crr_1985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => call_stmt_667_call_req_0); -- 
    ccr_2261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => call_stmt_778_call_req_1); -- 
    ccr_2275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => call_stmt_783_call_req_1); -- 
    cr_2321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => LOAD_next_pc1_795_load_0_req_1); -- 
    ccr_2289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => call_stmt_790_call_req_1); -- 
    req_2336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => MUX_883_inst_req_1); -- 
    ccr_2247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => call_stmt_771_call_req_1); -- 
    cr_2051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => STORE_next_pc1_675_store_0_req_1); -- 
    ccr_2065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => call_stmt_682_call_req_1); -- 
    ccr_2079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => call_stmt_688_call_req_1); -- 
    ccr_2093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => call_stmt_694_call_req_1); -- 
    ccr_2107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => call_stmt_701_call_req_1); -- 
    ccr_2121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => call_stmt_708_call_req_1); -- 
    ccr_2135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => call_stmt_715_call_req_1); -- 
    ccr_2149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => call_stmt_722_call_req_1); -- 
    ccr_2163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => call_stmt_729_call_req_1); -- 
    ccr_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => call_stmt_736_call_req_1); -- 
    ccr_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => call_stmt_743_call_req_1); -- 
    ccr_2205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => call_stmt_750_call_req_1); -- 
    ccr_2219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => call_stmt_757_call_req_1); -- 
    ccr_2233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(0), ack => call_stmt_764_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_667_sample_completed_
      -- CP-element group 1: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_667_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_667_Sample/cra
      -- 
    cra_1986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_667_call_ack_0, ack => try_CP_1972_elements(1)); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	48 
    -- CP-element group 2: 	51 
    -- CP-element group 2: 	69 
    -- CP-element group 2: 	54 
    -- CP-element group 2: 	56 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	21 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	27 
    -- CP-element group 2: 	30 
    -- CP-element group 2: 	33 
    -- CP-element group 2: 	36 
    -- CP-element group 2: 	39 
    -- CP-element group 2: 	42 
    -- CP-element group 2: 	45 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_667_update_completed_
      -- CP-element group 2: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_667_Update/$exit
      -- CP-element group 2: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_667_Update/cca
      -- CP-element group 2: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_783_sample_start_
      -- CP-element group 2: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_783_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_783_Sample/crr
      -- 
    cca_1991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_667_call_ack_1, ack => try_CP_1972_elements(2)); -- 
    crr_2270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(2), ack => call_stmt_783_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	69 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_672_sample_completed_
      -- CP-element group 3: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_672_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_672_Sample/cra
      -- 
    cra_2000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_672_call_ack_0, ack => try_CP_1972_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	48 
    -- CP-element group 4: 	51 
    -- CP-element group 4: 	70 
    -- CP-element group 4: 	56 
    -- CP-element group 4: 	15 
    -- CP-element group 4: 	18 
    -- CP-element group 4: 	21 
    -- CP-element group 4: 	24 
    -- CP-element group 4: 	27 
    -- CP-element group 4: 	30 
    -- CP-element group 4: 	33 
    -- CP-element group 4: 	36 
    -- CP-element group 4: 	39 
    -- CP-element group 4: 	42 
    -- CP-element group 4: 	45 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_672_update_completed_
      -- CP-element group 4: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_672_Update/$exit
      -- CP-element group 4: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_672_Update/cca
      -- 
    cca_2005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_672_call_ack_1, ack => try_CP_1972_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_676_sample_completed_
      -- CP-element group 5: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_676_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_676_Sample/cra
      -- 
    cra_2014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_676_call_ack_0, ack => try_CP_1972_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_676_update_completed_
      -- CP-element group 6: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_676_Update/$exit
      -- CP-element group 6: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_676_Update/cca
      -- 
    cca_2019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_676_call_ack_1, ack => try_CP_1972_elements(6)); -- 
    -- CP-element group 7:  join  transition  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (9) 
      -- CP-element group 7: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_sample_start_
      -- CP-element group 7: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_Sample/$entry
      -- CP-element group 7: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_Sample/STORE_next_pc1_675_Split/$entry
      -- CP-element group 7: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_Sample/STORE_next_pc1_675_Split/$exit
      -- CP-element group 7: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_Sample/STORE_next_pc1_675_Split/split_req
      -- CP-element group 7: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_Sample/STORE_next_pc1_675_Split/split_ack
      -- CP-element group 7: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_Sample/word_access_start/$entry
      -- CP-element group 7: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_Sample/word_access_start/word_0/$entry
      -- CP-element group 7: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_Sample/word_access_start/word_0/rr
      -- 
    rr_2040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(7), ack => STORE_next_pc1_675_store_0_req_0); -- 
    try_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 22) := "try_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try_CP_1972_elements(0) & try_CP_1972_elements(6);
      gj_try_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_1972_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	65 
    -- CP-element group 8:  members (5) 
      -- CP-element group 8: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_sample_completed_
      -- CP-element group 8: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_Sample/$exit
      -- CP-element group 8: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_Sample/word_access_start/$exit
      -- CP-element group 8: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_Sample/word_access_start/word_0/$exit
      -- CP-element group 8: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_Sample/word_access_start/word_0/ra
      -- 
    ra_2041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_next_pc1_675_store_0_ack_0, ack => try_CP_1972_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	83 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_update_completed_
      -- CP-element group 9: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_Update/$exit
      -- CP-element group 9: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_Update/word_access_complete/$exit
      -- CP-element group 9: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_Update/word_access_complete/word_0/$exit
      -- CP-element group 9: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_Update/word_access_complete/word_0/ca
      -- 
    ca_2052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_next_pc1_675_store_0_ack_1, ack => try_CP_1972_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	70 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_682_sample_completed_
      -- CP-element group 10: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_682_Sample/$exit
      -- CP-element group 10: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_682_Sample/cra
      -- 
    cra_2061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_682_call_ack_0, ack => try_CP_1972_elements(10)); -- 
    -- CP-element group 11:  fork  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	71 
    -- CP-element group 11: 	59 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_682_update_completed_
      -- CP-element group 11: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_682_Update/$exit
      -- CP-element group 11: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_682_Update/cca
      -- 
    cca_2066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_682_call_ack_1, ack => try_CP_1972_elements(11)); -- 
    -- CP-element group 12:  join  transition  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: 	71 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_688_sample_start_
      -- CP-element group 12: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_688_Sample/$entry
      -- CP-element group 12: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_688_Sample/crr
      -- 
    crr_2074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(12), ack => call_stmt_688_call_req_0); -- 
    try_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try_CP_1972_elements(2) & try_CP_1972_elements(71);
      gj_try_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_1972_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_688_sample_completed_
      -- CP-element group 13: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_688_Sample/$exit
      -- CP-element group 13: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_688_Sample/cra
      -- 
    cra_2075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_688_call_ack_0, ack => try_CP_1972_elements(13)); -- 
    -- CP-element group 14:  fork  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	0 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	68 
    -- CP-element group 14: 	72 
    -- CP-element group 14: 	59 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_688_update_completed_
      -- CP-element group 14: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_688_Update/$exit
      -- CP-element group 14: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_688_Update/cca
      -- 
    cca_2080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_688_call_ack_1, ack => try_CP_1972_elements(14)); -- 
    -- CP-element group 15:  join  transition  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: 	4 
    -- CP-element group 15: 	68 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_694_sample_start_
      -- CP-element group 15: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_694_Sample/$entry
      -- CP-element group 15: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_694_Sample/crr
      -- 
    crr_2088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(15), ack => call_stmt_694_call_req_0); -- 
    try_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try_CP_1972_elements(2) & try_CP_1972_elements(4) & try_CP_1972_elements(68);
      gj_try_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_1972_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_694_sample_completed_
      -- CP-element group 16: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_694_Sample/$exit
      -- CP-element group 16: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_694_Sample/cra
      -- 
    cra_2089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_694_call_ack_0, ack => try_CP_1972_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	59 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_694_update_completed_
      -- CP-element group 17: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_694_Update/$exit
      -- CP-element group 17: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_694_Update/cca
      -- 
    cca_2094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_694_call_ack_1, ack => try_CP_1972_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: 	4 
    -- CP-element group 18: 	72 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_701_sample_start_
      -- CP-element group 18: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_701_Sample/$entry
      -- CP-element group 18: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_701_Sample/crr
      -- 
    crr_2102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(18), ack => call_stmt_701_call_req_0); -- 
    try_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try_CP_1972_elements(2) & try_CP_1972_elements(4) & try_CP_1972_elements(72);
      gj_try_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_1972_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_701_sample_completed_
      -- CP-element group 19: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_701_Sample/$exit
      -- CP-element group 19: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_701_Sample/cra
      -- 
    cra_2103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_701_call_ack_0, ack => try_CP_1972_elements(19)); -- 
    -- CP-element group 20:  fork  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	73 
    -- CP-element group 20: 	59 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_701_update_completed_
      -- CP-element group 20: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_701_Update/$exit
      -- CP-element group 20: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_701_Update/cca
      -- 
    cca_2108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_701_call_ack_1, ack => try_CP_1972_elements(20)); -- 
    -- CP-element group 21:  join  transition  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	2 
    -- CP-element group 21: 	4 
    -- CP-element group 21: 	73 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_708_sample_start_
      -- CP-element group 21: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_708_Sample/$entry
      -- CP-element group 21: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_708_Sample/crr
      -- 
    crr_2116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(21), ack => call_stmt_708_call_req_0); -- 
    try_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try_CP_1972_elements(2) & try_CP_1972_elements(4) & try_CP_1972_elements(73);
      gj_try_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_1972_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_708_sample_completed_
      -- CP-element group 22: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_708_Sample/$exit
      -- CP-element group 22: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_708_Sample/cra
      -- 
    cra_2117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_708_call_ack_0, ack => try_CP_1972_elements(22)); -- 
    -- CP-element group 23:  fork  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	74 
    -- CP-element group 23: 	59 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_708_update_completed_
      -- CP-element group 23: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_708_Update/$exit
      -- CP-element group 23: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_708_Update/cca
      -- 
    cca_2122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_708_call_ack_1, ack => try_CP_1972_elements(23)); -- 
    -- CP-element group 24:  join  transition  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: 	4 
    -- CP-element group 24: 	74 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_715_sample_start_
      -- CP-element group 24: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_715_Sample/$entry
      -- CP-element group 24: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_715_Sample/crr
      -- 
    crr_2130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(24), ack => call_stmt_715_call_req_0); -- 
    try_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try_CP_1972_elements(2) & try_CP_1972_elements(4) & try_CP_1972_elements(74);
      gj_try_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_1972_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_715_sample_completed_
      -- CP-element group 25: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_715_Sample/$exit
      -- CP-element group 25: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_715_Sample/cra
      -- 
    cra_2131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_715_call_ack_0, ack => try_CP_1972_elements(25)); -- 
    -- CP-element group 26:  fork  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	0 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	75 
    -- CP-element group 26: 	59 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_715_update_completed_
      -- CP-element group 26: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_715_Update/$exit
      -- CP-element group 26: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_715_Update/cca
      -- 
    cca_2136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_715_call_ack_1, ack => try_CP_1972_elements(26)); -- 
    -- CP-element group 27:  join  transition  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: 	4 
    -- CP-element group 27: 	75 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_722_sample_start_
      -- CP-element group 27: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_722_Sample/$entry
      -- CP-element group 27: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_722_Sample/crr
      -- 
    crr_2144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(27), ack => call_stmt_722_call_req_0); -- 
    try_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try_CP_1972_elements(2) & try_CP_1972_elements(4) & try_CP_1972_elements(75);
      gj_try_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_1972_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_722_sample_completed_
      -- CP-element group 28: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_722_Sample/$exit
      -- CP-element group 28: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_722_Sample/cra
      -- 
    cra_2145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_722_call_ack_0, ack => try_CP_1972_elements(28)); -- 
    -- CP-element group 29:  fork  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	0 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	76 
    -- CP-element group 29: 	59 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_722_update_completed_
      -- CP-element group 29: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_722_Update/$exit
      -- CP-element group 29: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_722_Update/cca
      -- 
    cca_2150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_722_call_ack_1, ack => try_CP_1972_elements(29)); -- 
    -- CP-element group 30:  join  transition  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	2 
    -- CP-element group 30: 	4 
    -- CP-element group 30: 	76 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_729_sample_start_
      -- CP-element group 30: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_729_Sample/$entry
      -- CP-element group 30: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_729_Sample/crr
      -- 
    crr_2158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(30), ack => call_stmt_729_call_req_0); -- 
    try_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try_CP_1972_elements(2) & try_CP_1972_elements(4) & try_CP_1972_elements(76);
      gj_try_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_1972_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_729_sample_completed_
      -- CP-element group 31: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_729_Sample/$exit
      -- CP-element group 31: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_729_Sample/cra
      -- 
    cra_2159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_729_call_ack_0, ack => try_CP_1972_elements(31)); -- 
    -- CP-element group 32:  fork  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	77 
    -- CP-element group 32: 	59 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_729_update_completed_
      -- CP-element group 32: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_729_Update/$exit
      -- CP-element group 32: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_729_Update/cca
      -- 
    cca_2164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_729_call_ack_1, ack => try_CP_1972_elements(32)); -- 
    -- CP-element group 33:  join  transition  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	2 
    -- CP-element group 33: 	4 
    -- CP-element group 33: 	77 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_736_sample_start_
      -- CP-element group 33: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_736_Sample/$entry
      -- CP-element group 33: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_736_Sample/crr
      -- 
    crr_2172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(33), ack => call_stmt_736_call_req_0); -- 
    try_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try_CP_1972_elements(2) & try_CP_1972_elements(4) & try_CP_1972_elements(77);
      gj_try_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_1972_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_736_sample_completed_
      -- CP-element group 34: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_736_Sample/$exit
      -- CP-element group 34: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_736_Sample/cra
      -- 
    cra_2173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_736_call_ack_0, ack => try_CP_1972_elements(34)); -- 
    -- CP-element group 35:  fork  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	0 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	78 
    -- CP-element group 35: 	59 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_736_update_completed_
      -- CP-element group 35: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_736_Update/$exit
      -- CP-element group 35: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_736_Update/cca
      -- 
    cca_2178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_736_call_ack_1, ack => try_CP_1972_elements(35)); -- 
    -- CP-element group 36:  join  transition  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	2 
    -- CP-element group 36: 	4 
    -- CP-element group 36: 	78 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_743_sample_start_
      -- CP-element group 36: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_743_Sample/$entry
      -- CP-element group 36: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_743_Sample/crr
      -- 
    crr_2186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(36), ack => call_stmt_743_call_req_0); -- 
    try_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try_CP_1972_elements(2) & try_CP_1972_elements(4) & try_CP_1972_elements(78);
      gj_try_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_1972_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_743_sample_completed_
      -- CP-element group 37: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_743_Sample/$exit
      -- CP-element group 37: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_743_Sample/cra
      -- 
    cra_2187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_743_call_ack_0, ack => try_CP_1972_elements(37)); -- 
    -- CP-element group 38:  fork  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	0 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	79 
    -- CP-element group 38: 	59 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_743_update_completed_
      -- CP-element group 38: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_743_Update/$exit
      -- CP-element group 38: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_743_Update/cca
      -- 
    cca_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_743_call_ack_1, ack => try_CP_1972_elements(38)); -- 
    -- CP-element group 39:  join  transition  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	2 
    -- CP-element group 39: 	4 
    -- CP-element group 39: 	79 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_750_sample_start_
      -- CP-element group 39: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_750_Sample/$entry
      -- CP-element group 39: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_750_Sample/crr
      -- 
    crr_2200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(39), ack => call_stmt_750_call_req_0); -- 
    try_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try_CP_1972_elements(2) & try_CP_1972_elements(4) & try_CP_1972_elements(79);
      gj_try_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_1972_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_750_sample_completed_
      -- CP-element group 40: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_750_Sample/$exit
      -- CP-element group 40: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_750_Sample/cra
      -- 
    cra_2201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_750_call_ack_0, ack => try_CP_1972_elements(40)); -- 
    -- CP-element group 41:  fork  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	0 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	80 
    -- CP-element group 41: 	59 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_750_update_completed_
      -- CP-element group 41: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_750_Update/$exit
      -- CP-element group 41: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_750_Update/cca
      -- 
    cca_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_750_call_ack_1, ack => try_CP_1972_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	2 
    -- CP-element group 42: 	4 
    -- CP-element group 42: 	80 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_757_sample_start_
      -- CP-element group 42: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_757_Sample/$entry
      -- CP-element group 42: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_757_Sample/crr
      -- 
    crr_2214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(42), ack => call_stmt_757_call_req_0); -- 
    try_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try_CP_1972_elements(2) & try_CP_1972_elements(4) & try_CP_1972_elements(80);
      gj_try_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_1972_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_757_sample_completed_
      -- CP-element group 43: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_757_Sample/$exit
      -- CP-element group 43: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_757_Sample/cra
      -- 
    cra_2215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_757_call_ack_0, ack => try_CP_1972_elements(43)); -- 
    -- CP-element group 44:  fork  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	81 
    -- CP-element group 44: 	59 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_757_update_completed_
      -- CP-element group 44: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_757_Update/$exit
      -- CP-element group 44: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_757_Update/cca
      -- 
    cca_2220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_757_call_ack_1, ack => try_CP_1972_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	2 
    -- CP-element group 45: 	4 
    -- CP-element group 45: 	65 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_764_sample_start_
      -- CP-element group 45: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_764_Sample/$entry
      -- CP-element group 45: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_764_Sample/crr
      -- 
    crr_2228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(45), ack => call_stmt_764_call_req_0); -- 
    try_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try_CP_1972_elements(2) & try_CP_1972_elements(4) & try_CP_1972_elements(65);
      gj_try_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_1972_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_764_sample_completed_
      -- CP-element group 46: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_764_Sample/$exit
      -- CP-element group 46: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_764_Sample/cra
      -- 
    cra_2229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_764_call_ack_0, ack => try_CP_1972_elements(46)); -- 
    -- CP-element group 47:  fork  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	0 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	66 
    -- CP-element group 47: 	59 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_764_update_completed_
      -- CP-element group 47: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_764_Update/$exit
      -- CP-element group 47: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_764_Update/cca
      -- 
    cca_2234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_764_call_ack_1, ack => try_CP_1972_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	2 
    -- CP-element group 48: 	4 
    -- CP-element group 48: 	66 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_771_sample_start_
      -- CP-element group 48: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_771_Sample/$entry
      -- CP-element group 48: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_771_Sample/crr
      -- 
    crr_2242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(48), ack => call_stmt_771_call_req_0); -- 
    try_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try_CP_1972_elements(2) & try_CP_1972_elements(4) & try_CP_1972_elements(66);
      gj_try_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_1972_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_771_sample_completed_
      -- CP-element group 49: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_771_Sample/$exit
      -- CP-element group 49: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_771_Sample/cra
      -- 
    cra_2243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_771_call_ack_0, ack => try_CP_1972_elements(49)); -- 
    -- CP-element group 50:  fork  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	0 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	67 
    -- CP-element group 50: 	59 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_771_update_completed_
      -- CP-element group 50: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_771_Update/$exit
      -- CP-element group 50: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_771_Update/cca
      -- 
    cca_2248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_771_call_ack_1, ack => try_CP_1972_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	2 
    -- CP-element group 51: 	4 
    -- CP-element group 51: 	81 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_778_sample_start_
      -- CP-element group 51: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_778_Sample/$entry
      -- CP-element group 51: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_778_Sample/crr
      -- 
    crr_2256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(51), ack => call_stmt_778_call_req_0); -- 
    try_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try_CP_1972_elements(2) & try_CP_1972_elements(4) & try_CP_1972_elements(81);
      gj_try_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_1972_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_778_sample_completed_
      -- CP-element group 52: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_778_Sample/$exit
      -- CP-element group 52: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_778_Sample/cra
      -- 
    cra_2257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_778_call_ack_0, ack => try_CP_1972_elements(52)); -- 
    -- CP-element group 53:  fork  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	0 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	82 
    -- CP-element group 53: 	59 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_778_update_completed_
      -- CP-element group 53: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_778_Update/$exit
      -- CP-element group 53: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_778_Update/cca
      -- 
    cca_2262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_778_call_ack_1, ack => try_CP_1972_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	2 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_783_sample_completed_
      -- CP-element group 54: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_783_Sample/$exit
      -- CP-element group 54: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_783_Sample/cra
      -- 
    cra_2271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_783_call_ack_0, ack => try_CP_1972_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	0 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	59 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_783_update_completed_
      -- CP-element group 55: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_783_Update/$exit
      -- CP-element group 55: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_783_Update/cca
      -- 
    cca_2276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_783_call_ack_1, ack => try_CP_1972_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	2 
    -- CP-element group 56: 	4 
    -- CP-element group 56: 	82 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_790_sample_start_
      -- CP-element group 56: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_790_Sample/$entry
      -- CP-element group 56: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_790_Sample/crr
      -- 
    crr_2284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(56), ack => call_stmt_790_call_req_0); -- 
    try_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= try_CP_1972_elements(2) & try_CP_1972_elements(4) & try_CP_1972_elements(82);
      gj_try_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_1972_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_790_sample_completed_
      -- CP-element group 57: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_790_Sample/$exit
      -- CP-element group 57: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_790_Sample/cra
      -- 
    cra_2285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_790_call_ack_0, ack => try_CP_1972_elements(57)); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	0 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_790_update_completed_
      -- CP-element group 58: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_790_Update/$exit
      -- CP-element group 58: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_790_Update/cca
      -- 
    cca_2290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_790_call_ack_1, ack => try_CP_1972_elements(58)); -- 
    -- CP-element group 59:  join  transition  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	50 
    -- CP-element group 59: 	47 
    -- CP-element group 59: 	53 
    -- CP-element group 59: 	58 
    -- CP-element group 59: 	55 
    -- CP-element group 59: 	62 
    -- CP-element group 59: 	11 
    -- CP-element group 59: 	14 
    -- CP-element group 59: 	17 
    -- CP-element group 59: 	20 
    -- CP-element group 59: 	23 
    -- CP-element group 59: 	26 
    -- CP-element group 59: 	29 
    -- CP-element group 59: 	32 
    -- CP-element group 59: 	35 
    -- CP-element group 59: 	38 
    -- CP-element group 59: 	41 
    -- CP-element group 59: 	44 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	63 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 assign_stmt_560_to_assign_stmt_884/MUX_883_sample_start_
      -- CP-element group 59: 	 assign_stmt_560_to_assign_stmt_884/MUX_883_start/req
      -- CP-element group 59: 	 assign_stmt_560_to_assign_stmt_884/MUX_883_start/$entry
      -- 
    req_2331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(59), ack => MUX_883_inst_req_0); -- 
    try_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 17) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1);
      constant place_markings: IntegerArray(0 to 17)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0);
      constant place_delays: IntegerArray(0 to 17) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 18); -- 
    begin -- 
      preds <= try_CP_1972_elements(50) & try_CP_1972_elements(47) & try_CP_1972_elements(53) & try_CP_1972_elements(58) & try_CP_1972_elements(55) & try_CP_1972_elements(62) & try_CP_1972_elements(11) & try_CP_1972_elements(14) & try_CP_1972_elements(17) & try_CP_1972_elements(20) & try_CP_1972_elements(23) & try_CP_1972_elements(26) & try_CP_1972_elements(29) & try_CP_1972_elements(32) & try_CP_1972_elements(35) & try_CP_1972_elements(38) & try_CP_1972_elements(41) & try_CP_1972_elements(44);
      gj_try_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 18, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_1972_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  join  transition  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: 	67 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (5) 
      -- CP-element group 60: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_Sample/word_access_start/word_0/rr
      -- CP-element group 60: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_Sample/word_access_start/word_0/$entry
      -- CP-element group 60: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_sample_start_
      -- CP-element group 60: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_Sample/word_access_start/$entry
      -- CP-element group 60: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_Sample/$entry
      -- 
    rr_2310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(60), ack => LOAD_next_pc1_795_load_0_req_0); -- 
    try_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try_CP_1972_elements(0) & try_CP_1972_elements(67);
      gj_try_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_1972_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (5) 
      -- CP-element group 61: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_Sample/$exit
      -- CP-element group 61: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_Sample/word_access_start/word_0/$exit
      -- CP-element group 61: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_sample_completed_
      -- CP-element group 61: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_Sample/word_access_start/word_0/ra
      -- CP-element group 61: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_Sample/word_access_start/$exit
      -- 
    ra_2311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_next_pc1_795_load_0_ack_0, ack => try_CP_1972_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	0 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	59 
    -- CP-element group 62:  members (9) 
      -- CP-element group 62: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_Update/word_access_complete/word_0/$exit
      -- CP-element group 62: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_Update/word_access_complete/word_0/ca
      -- CP-element group 62: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_Update/LOAD_next_pc1_795_Merge/$entry
      -- CP-element group 62: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_Update/$exit
      -- CP-element group 62: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_Update/LOAD_next_pc1_795_Merge/$exit
      -- CP-element group 62: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_Update/LOAD_next_pc1_795_Merge/merge_req
      -- CP-element group 62: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_Update/LOAD_next_pc1_795_Merge/merge_ack
      -- CP-element group 62: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_Update/word_access_complete/$exit
      -- CP-element group 62: 	 assign_stmt_560_to_assign_stmt_884/LOAD_next_pc1_795_update_completed_
      -- 
    ca_2322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_next_pc1_795_load_0_ack_1, ack => try_CP_1972_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	59 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 assign_stmt_560_to_assign_stmt_884/MUX_883_sample_completed_
      -- CP-element group 63: 	 assign_stmt_560_to_assign_stmt_884/MUX_883_start/ack
      -- CP-element group 63: 	 assign_stmt_560_to_assign_stmt_884/MUX_883_start/$exit
      -- 
    ack_2332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_883_inst_ack_0, ack => try_CP_1972_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	0 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	83 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 assign_stmt_560_to_assign_stmt_884/MUX_883_update_completed_
      -- CP-element group 64: 	 assign_stmt_560_to_assign_stmt_884/MUX_883_complete/ack
      -- CP-element group 64: 	 assign_stmt_560_to_assign_stmt_884/MUX_883_complete/$exit
      -- 
    ack_2337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_883_inst_ack_1, ack => try_CP_1972_elements(64)); -- 
    -- CP-element group 65:  transition  delay-element  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	8 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	45 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 assign_stmt_560_to_assign_stmt_884/STORE_next_pc1_675_call_stmt_764_delay
      -- 
    -- Element group try_CP_1972_elements(65) is a control-delay.
    cp_element_65_delay: control_delay_element  generic map(name => " 65_delay", delay_value => 1)  port map(req => try_CP_1972_elements(8), ack => try_CP_1972_elements(65), clk => clk, reset =>reset);
    -- CP-element group 66:  transition  delay-element  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	47 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	48 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_764_call_stmt_771_delay
      -- 
    -- Element group try_CP_1972_elements(66) is a control-delay.
    cp_element_66_delay: control_delay_element  generic map(name => " 66_delay", delay_value => 1)  port map(req => try_CP_1972_elements(47), ack => try_CP_1972_elements(66), clk => clk, reset =>reset);
    -- CP-element group 67:  transition  delay-element  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	50 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	60 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_771_LOAD_next_pc1_795_delay
      -- 
    -- Element group try_CP_1972_elements(67) is a control-delay.
    cp_element_67_delay: control_delay_element  generic map(name => " 67_delay", delay_value => 1)  port map(req => try_CP_1972_elements(50), ack => try_CP_1972_elements(67), clk => clk, reset =>reset);
    -- CP-element group 68:  transition  delay-element  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	14 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	15 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_688_call_stmt_694_delay
      -- 
    -- Element group try_CP_1972_elements(68) is a control-delay.
    cp_element_68_delay: control_delay_element  generic map(name => " 68_delay", delay_value => 1)  port map(req => try_CP_1972_elements(14), ack => try_CP_1972_elements(68), clk => clk, reset =>reset);
    -- CP-element group 69:  transition  output  delay-element  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	2 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	3 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_672_sample_start_
      -- CP-element group 69: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_672_Sample/$entry
      -- CP-element group 69: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_672_Sample/crr
      -- CP-element group 69: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_667_call_stmt_672_delay
      -- 
    crr_1999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(69), ack => call_stmt_672_call_req_0); -- 
    -- Element group try_CP_1972_elements(69) is a control-delay.
    cp_element_69_delay: control_delay_element  generic map(name => " 69_delay", delay_value => 1)  port map(req => try_CP_1972_elements(2), ack => try_CP_1972_elements(69), clk => clk, reset =>reset);
    -- CP-element group 70:  transition  output  delay-element  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	4 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	10 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_682_sample_start_
      -- CP-element group 70: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_682_Sample/$entry
      -- CP-element group 70: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_682_Sample/crr
      -- CP-element group 70: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_672_call_stmt_682_delay
      -- 
    crr_2060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try_CP_1972_elements(70), ack => call_stmt_682_call_req_0); -- 
    -- Element group try_CP_1972_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => try_CP_1972_elements(4), ack => try_CP_1972_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  transition  delay-element  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	11 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	12 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_682_call_stmt_688_delay
      -- 
    -- Element group try_CP_1972_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => try_CP_1972_elements(11), ack => try_CP_1972_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  transition  delay-element  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	14 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	18 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_688_call_stmt_701_delay
      -- 
    -- Element group try_CP_1972_elements(72) is a control-delay.
    cp_element_72_delay: control_delay_element  generic map(name => " 72_delay", delay_value => 1)  port map(req => try_CP_1972_elements(14), ack => try_CP_1972_elements(72), clk => clk, reset =>reset);
    -- CP-element group 73:  transition  delay-element  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	20 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	21 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_701_call_stmt_708_delay
      -- 
    -- Element group try_CP_1972_elements(73) is a control-delay.
    cp_element_73_delay: control_delay_element  generic map(name => " 73_delay", delay_value => 1)  port map(req => try_CP_1972_elements(20), ack => try_CP_1972_elements(73), clk => clk, reset =>reset);
    -- CP-element group 74:  transition  delay-element  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	23 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	24 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_708_call_stmt_715_delay
      -- 
    -- Element group try_CP_1972_elements(74) is a control-delay.
    cp_element_74_delay: control_delay_element  generic map(name => " 74_delay", delay_value => 1)  port map(req => try_CP_1972_elements(23), ack => try_CP_1972_elements(74), clk => clk, reset =>reset);
    -- CP-element group 75:  transition  delay-element  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	26 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	27 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_715_call_stmt_722_delay
      -- 
    -- Element group try_CP_1972_elements(75) is a control-delay.
    cp_element_75_delay: control_delay_element  generic map(name => " 75_delay", delay_value => 1)  port map(req => try_CP_1972_elements(26), ack => try_CP_1972_elements(75), clk => clk, reset =>reset);
    -- CP-element group 76:  transition  delay-element  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	29 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	30 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_722_call_stmt_729_delay
      -- 
    -- Element group try_CP_1972_elements(76) is a control-delay.
    cp_element_76_delay: control_delay_element  generic map(name => " 76_delay", delay_value => 1)  port map(req => try_CP_1972_elements(29), ack => try_CP_1972_elements(76), clk => clk, reset =>reset);
    -- CP-element group 77:  transition  delay-element  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	32 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	33 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_729_call_stmt_736_delay
      -- 
    -- Element group try_CP_1972_elements(77) is a control-delay.
    cp_element_77_delay: control_delay_element  generic map(name => " 77_delay", delay_value => 1)  port map(req => try_CP_1972_elements(32), ack => try_CP_1972_elements(77), clk => clk, reset =>reset);
    -- CP-element group 78:  transition  delay-element  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	35 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	36 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_736_call_stmt_743_delay
      -- 
    -- Element group try_CP_1972_elements(78) is a control-delay.
    cp_element_78_delay: control_delay_element  generic map(name => " 78_delay", delay_value => 1)  port map(req => try_CP_1972_elements(35), ack => try_CP_1972_elements(78), clk => clk, reset =>reset);
    -- CP-element group 79:  transition  delay-element  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	38 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	39 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_743_call_stmt_750_delay
      -- 
    -- Element group try_CP_1972_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => try_CP_1972_elements(38), ack => try_CP_1972_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  transition  delay-element  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	41 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	42 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_750_call_stmt_757_delay
      -- 
    -- Element group try_CP_1972_elements(80) is a control-delay.
    cp_element_80_delay: control_delay_element  generic map(name => " 80_delay", delay_value => 1)  port map(req => try_CP_1972_elements(41), ack => try_CP_1972_elements(80), clk => clk, reset =>reset);
    -- CP-element group 81:  transition  delay-element  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	44 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	51 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_757_call_stmt_778_delay
      -- 
    -- Element group try_CP_1972_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => try_CP_1972_elements(44), ack => try_CP_1972_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  transition  delay-element  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	53 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	56 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 assign_stmt_560_to_assign_stmt_884/call_stmt_778_call_stmt_790_delay
      -- 
    -- Element group try_CP_1972_elements(82) is a control-delay.
    cp_element_82_delay: control_delay_element  generic map(name => " 82_delay", delay_value => 1)  port map(req => try_CP_1972_elements(53), ack => try_CP_1972_elements(82), clk => clk, reset =>reset);
    -- CP-element group 83:  join  transition  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	64 
    -- CP-element group 83: 	9 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 $exit
      -- CP-element group 83: 	 assign_stmt_560_to_assign_stmt_884/$exit
      -- 
    try_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 23) := "try_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try_CP_1972_elements(64) & try_CP_1972_elements(9);
      gj_try_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try_CP_1972_elements(83), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u8_u1_794_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_798_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_802_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_806_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_810_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_814_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_818_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_822_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_826_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_830_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_834_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_838_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_842_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_846_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_850_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_854_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_858_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_862_wire : std_logic_vector(0 downto 0);
    signal LOAD_next_pc1_795_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_next_pc1_795_wire : std_logic_vector(7 downto 0);
    signal LOAD_next_pc1_795_word_address_0 : std_logic_vector(0 downto 0);
    signal MUX_866_wire : std_logic_vector(7 downto 0);
    signal MUX_867_wire : std_logic_vector(7 downto 0);
    signal MUX_868_wire : std_logic_vector(7 downto 0);
    signal MUX_869_wire : std_logic_vector(7 downto 0);
    signal MUX_870_wire : std_logic_vector(7 downto 0);
    signal MUX_871_wire : std_logic_vector(7 downto 0);
    signal MUX_872_wire : std_logic_vector(7 downto 0);
    signal MUX_873_wire : std_logic_vector(7 downto 0);
    signal MUX_874_wire : std_logic_vector(7 downto 0);
    signal MUX_875_wire : std_logic_vector(7 downto 0);
    signal MUX_876_wire : std_logic_vector(7 downto 0);
    signal MUX_877_wire : std_logic_vector(7 downto 0);
    signal MUX_878_wire : std_logic_vector(7 downto 0);
    signal MUX_879_wire : std_logic_vector(7 downto 0);
    signal MUX_880_wire : std_logic_vector(7 downto 0);
    signal MUX_881_wire : std_logic_vector(7 downto 0);
    signal MUX_882_wire : std_logic_vector(7 downto 0);
    signal STORE_next_pc1_675_data_0 : std_logic_vector(7 downto 0);
    signal STORE_next_pc1_675_wire : std_logic_vector(7 downto 0);
    signal STORE_next_pc1_675_word_address_0 : std_logic_vector(0 downto 0);
    signal add1_617 : std_logic_vector(0 downto 0);
    signal and1_597 : std_logic_vector(0 downto 0);
    signal bn1_647 : std_logic_vector(0 downto 0);
    signal bz1_642 : std_logic_vector(0 downto 0);
    signal call1_652 : std_logic_vector(0 downto 0);
    signal cmp1_662 : std_logic_vector(0 downto 0);
    signal halt1_577 : std_logic_vector(0 downto 0);
    signal jmp1_657 : std_logic_vector(0 downto 0);
    signal konst_575_wire_constant : std_logic_vector(7 downto 0);
    signal konst_580_wire_constant : std_logic_vector(7 downto 0);
    signal konst_585_wire_constant : std_logic_vector(7 downto 0);
    signal konst_590_wire_constant : std_logic_vector(7 downto 0);
    signal konst_595_wire_constant : std_logic_vector(7 downto 0);
    signal konst_600_wire_constant : std_logic_vector(7 downto 0);
    signal konst_605_wire_constant : std_logic_vector(7 downto 0);
    signal konst_610_wire_constant : std_logic_vector(7 downto 0);
    signal konst_615_wire_constant : std_logic_vector(7 downto 0);
    signal konst_620_wire_constant : std_logic_vector(7 downto 0);
    signal konst_625_wire_constant : std_logic_vector(7 downto 0);
    signal konst_630_wire_constant : std_logic_vector(7 downto 0);
    signal konst_635_wire_constant : std_logic_vector(7 downto 0);
    signal konst_640_wire_constant : std_logic_vector(7 downto 0);
    signal konst_645_wire_constant : std_logic_vector(7 downto 0);
    signal konst_650_wire_constant : std_logic_vector(7 downto 0);
    signal konst_655_wire_constant : std_logic_vector(7 downto 0);
    signal konst_660_wire_constant : std_logic_vector(7 downto 0);
    signal konst_663_wire_constant : std_logic_vector(0 downto 0);
    signal konst_665_wire_constant : std_logic_vector(31 downto 0);
    signal konst_668_wire_constant : std_logic_vector(0 downto 0);
    signal konst_670_wire_constant : std_logic_vector(31 downto 0);
    signal konst_793_wire_constant : std_logic_vector(7 downto 0);
    signal konst_797_wire_constant : std_logic_vector(7 downto 0);
    signal konst_801_wire_constant : std_logic_vector(7 downto 0);
    signal konst_805_wire_constant : std_logic_vector(7 downto 0);
    signal konst_809_wire_constant : std_logic_vector(7 downto 0);
    signal konst_813_wire_constant : std_logic_vector(7 downto 0);
    signal konst_817_wire_constant : std_logic_vector(7 downto 0);
    signal konst_821_wire_constant : std_logic_vector(7 downto 0);
    signal konst_825_wire_constant : std_logic_vector(7 downto 0);
    signal konst_829_wire_constant : std_logic_vector(7 downto 0);
    signal konst_833_wire_constant : std_logic_vector(7 downto 0);
    signal konst_837_wire_constant : std_logic_vector(7 downto 0);
    signal konst_841_wire_constant : std_logic_vector(7 downto 0);
    signal konst_845_wire_constant : std_logic_vector(7 downto 0);
    signal konst_849_wire_constant : std_logic_vector(7 downto 0);
    signal konst_853_wire_constant : std_logic_vector(7 downto 0);
    signal konst_857_wire_constant : std_logic_vector(7 downto 0);
    signal konst_861_wire_constant : std_logic_vector(7 downto 0);
    signal load1_587 : std_logic_vector(0 downto 0);
    signal next_pc10_736 : std_logic_vector(7 downto 0);
    signal next_pc11_743 : std_logic_vector(7 downto 0);
    signal next_pc12_750 : std_logic_vector(7 downto 0);
    signal next_pc13_757 : std_logic_vector(7 downto 0);
    signal next_pc14_764 : std_logic_vector(7 downto 0);
    signal next_pc15_771 : std_logic_vector(7 downto 0);
    signal next_pc16_778 : std_logic_vector(7 downto 0);
    signal next_pc17_783 : std_logic_vector(7 downto 0);
    signal next_pc18_790 : std_logic_vector(7 downto 0);
    signal next_pc2_682 : std_logic_vector(7 downto 0);
    signal next_pc3_688 : std_logic_vector(7 downto 0);
    signal next_pc4_694 : std_logic_vector(7 downto 0);
    signal next_pc5_701 : std_logic_vector(7 downto 0);
    signal next_pc6_708 : std_logic_vector(7 downto 0);
    signal next_pc7_715 : std_logic_vector(7 downto 0);
    signal next_pc8_722 : std_logic_vector(7 downto 0);
    signal next_pc9_729 : std_logic_vector(7 downto 0);
    signal op_560 : std_logic_vector(7 downto 0);
    signal or1_602 : std_logic_vector(0 downto 0);
    signal rd_572 : std_logic_vector(7 downto 0);
    signal rs1_564 : std_logic_vector(7 downto 0);
    signal rs1_data_667 : std_logic_vector(31 downto 0);
    signal rs2_568 : std_logic_vector(7 downto 0);
    signal rs2_data_672 : std_logic_vector(31 downto 0);
    signal sbir1_582 : std_logic_vector(0 downto 0);
    signal sll1_627 : std_logic_vector(0 downto 0);
    signal sra1_637 : std_logic_vector(0 downto 0);
    signal srl1_632 : std_logic_vector(0 downto 0);
    signal store1_592 : std_logic_vector(0 downto 0);
    signal sub1_622 : std_logic_vector(0 downto 0);
    signal type_cast_865_wire_constant : std_logic_vector(7 downto 0);
    signal xnor1_607 : std_logic_vector(0 downto 0);
    signal xor1_612 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_next_pc1_795_word_address_0 <= "0";
    STORE_next_pc1_675_word_address_0 <= "0";
    konst_575_wire_constant <= "00000001";
    konst_580_wire_constant <= "00000010";
    konst_585_wire_constant <= "00000011";
    konst_590_wire_constant <= "00000100";
    konst_595_wire_constant <= "00000101";
    konst_600_wire_constant <= "00000110";
    konst_605_wire_constant <= "00000111";
    konst_610_wire_constant <= "00001000";
    konst_615_wire_constant <= "00001001";
    konst_620_wire_constant <= "00001010";
    konst_625_wire_constant <= "00001011";
    konst_630_wire_constant <= "00001100";
    konst_635_wire_constant <= "00001101";
    konst_640_wire_constant <= "00001110";
    konst_645_wire_constant <= "00001111";
    konst_650_wire_constant <= "00010000";
    konst_655_wire_constant <= "00010001";
    konst_660_wire_constant <= "00010010";
    konst_663_wire_constant <= "1";
    konst_665_wire_constant <= "00000000000000000000000000000000";
    konst_668_wire_constant <= "1";
    konst_670_wire_constant <= "00000000000000000000000000000000";
    konst_793_wire_constant <= "00000001";
    konst_797_wire_constant <= "00000010";
    konst_801_wire_constant <= "00000011";
    konst_805_wire_constant <= "00000100";
    konst_809_wire_constant <= "00000101";
    konst_813_wire_constant <= "00000110";
    konst_817_wire_constant <= "00000111";
    konst_821_wire_constant <= "00001000";
    konst_825_wire_constant <= "00001001";
    konst_829_wire_constant <= "00001010";
    konst_833_wire_constant <= "00001011";
    konst_837_wire_constant <= "00001100";
    konst_841_wire_constant <= "00001101";
    konst_845_wire_constant <= "00001110";
    konst_849_wire_constant <= "00001111";
    konst_853_wire_constant <= "00010000";
    konst_857_wire_constant <= "00010001";
    konst_861_wire_constant <= "00010010";
    type_cast_865_wire_constant <= "00000000";
    -- flow-through select operator MUX_866_inst
    MUX_866_wire <= next_pc18_790 when (EQ_u8_u1_862_wire(0) /=  '0') else type_cast_865_wire_constant;
    -- flow-through select operator MUX_867_inst
    MUX_867_wire <= next_pc17_783 when (EQ_u8_u1_858_wire(0) /=  '0') else MUX_866_wire;
    -- flow-through select operator MUX_868_inst
    MUX_868_wire <= next_pc16_778 when (EQ_u8_u1_854_wire(0) /=  '0') else MUX_867_wire;
    -- flow-through select operator MUX_869_inst
    MUX_869_wire <= next_pc15_771 when (EQ_u8_u1_850_wire(0) /=  '0') else MUX_868_wire;
    -- flow-through select operator MUX_870_inst
    MUX_870_wire <= next_pc14_764 when (EQ_u8_u1_846_wire(0) /=  '0') else MUX_869_wire;
    -- flow-through select operator MUX_871_inst
    MUX_871_wire <= next_pc13_757 when (EQ_u8_u1_842_wire(0) /=  '0') else MUX_870_wire;
    -- flow-through select operator MUX_872_inst
    MUX_872_wire <= next_pc12_750 when (EQ_u8_u1_838_wire(0) /=  '0') else MUX_871_wire;
    -- flow-through select operator MUX_873_inst
    MUX_873_wire <= next_pc11_743 when (EQ_u8_u1_834_wire(0) /=  '0') else MUX_872_wire;
    -- flow-through select operator MUX_874_inst
    MUX_874_wire <= next_pc10_736 when (EQ_u8_u1_830_wire(0) /=  '0') else MUX_873_wire;
    -- flow-through select operator MUX_875_inst
    MUX_875_wire <= next_pc9_729 when (EQ_u8_u1_826_wire(0) /=  '0') else MUX_874_wire;
    -- flow-through select operator MUX_876_inst
    MUX_876_wire <= next_pc8_722 when (EQ_u8_u1_822_wire(0) /=  '0') else MUX_875_wire;
    -- flow-through select operator MUX_877_inst
    MUX_877_wire <= next_pc7_715 when (EQ_u8_u1_818_wire(0) /=  '0') else MUX_876_wire;
    -- flow-through select operator MUX_878_inst
    MUX_878_wire <= next_pc6_708 when (EQ_u8_u1_814_wire(0) /=  '0') else MUX_877_wire;
    -- flow-through select operator MUX_879_inst
    MUX_879_wire <= next_pc5_701 when (EQ_u8_u1_810_wire(0) /=  '0') else MUX_878_wire;
    -- flow-through select operator MUX_880_inst
    MUX_880_wire <= next_pc4_694 when (EQ_u8_u1_806_wire(0) /=  '0') else MUX_879_wire;
    -- flow-through select operator MUX_881_inst
    MUX_881_wire <= next_pc3_688 when (EQ_u8_u1_802_wire(0) /=  '0') else MUX_880_wire;
    -- flow-through select operator MUX_882_inst
    MUX_882_wire <= next_pc2_682 when (EQ_u8_u1_798_wire(0) /=  '0') else MUX_881_wire;
    MUX_883_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_883_inst_req_0;
      MUX_883_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_883_inst_req_1;
      MUX_883_inst_ack_1<= update_ack(0);
      MUX_883_inst: SelectSplitProtocol generic map(name => "MUX_883_inst", data_width => 8, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => LOAD_next_pc1_795_wire, y => MUX_882_wire, sel => EQ_u8_u1_794_wire, z => next_pc_buffer, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through slice operator slice_559_inst
    op_560 <= inst_buffer(31 downto 24);
    -- flow-through slice operator slice_563_inst
    rs1_564 <= inst_buffer(23 downto 16);
    -- flow-through slice operator slice_567_inst
    rs2_568 <= inst_buffer(15 downto 8);
    -- flow-through slice operator slice_571_inst
    rd_572 <= inst_buffer(7 downto 0);
    -- equivalence LOAD_next_pc1_795_gather_scatter
    process(LOAD_next_pc1_795_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_next_pc1_795_data_0;
      ov(7 downto 0) := iv;
      LOAD_next_pc1_795_wire <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_next_pc1_675_gather_scatter
    process(STORE_next_pc1_675_wire) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := STORE_next_pc1_675_wire;
      ov(7 downto 0) := iv;
      STORE_next_pc1_675_data_0 <= ov(7 downto 0);
      --
    end process;
    -- binary operator EQ_u8_u1_576_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_575_wire_constant, tmp_var);
      halt1_577 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_581_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_580_wire_constant, tmp_var);
      sbir1_582 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_586_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_585_wire_constant, tmp_var);
      load1_587 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_591_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_590_wire_constant, tmp_var);
      store1_592 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_596_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_595_wire_constant, tmp_var);
      and1_597 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_601_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_600_wire_constant, tmp_var);
      or1_602 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_606_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_605_wire_constant, tmp_var);
      xnor1_607 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_611_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_610_wire_constant, tmp_var);
      xor1_612 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_616_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_615_wire_constant, tmp_var);
      add1_617 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_621_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_620_wire_constant, tmp_var);
      sub1_622 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_626_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_625_wire_constant, tmp_var);
      sll1_627 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_631_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_630_wire_constant, tmp_var);
      srl1_632 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_636_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_635_wire_constant, tmp_var);
      sra1_637 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_641_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_640_wire_constant, tmp_var);
      bz1_642 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_646_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_645_wire_constant, tmp_var);
      bn1_647 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_651_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_650_wire_constant, tmp_var);
      call1_652 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_656_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_655_wire_constant, tmp_var);
      jmp1_657 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_661_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_660_wire_constant, tmp_var);
      cmp1_662 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_794_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_793_wire_constant, tmp_var);
      EQ_u8_u1_794_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_798_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_797_wire_constant, tmp_var);
      EQ_u8_u1_798_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_802_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_801_wire_constant, tmp_var);
      EQ_u8_u1_802_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_806_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_805_wire_constant, tmp_var);
      EQ_u8_u1_806_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_810_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_809_wire_constant, tmp_var);
      EQ_u8_u1_810_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_814_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_813_wire_constant, tmp_var);
      EQ_u8_u1_814_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_818_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_817_wire_constant, tmp_var);
      EQ_u8_u1_818_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_822_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_821_wire_constant, tmp_var);
      EQ_u8_u1_822_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_826_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_825_wire_constant, tmp_var);
      EQ_u8_u1_826_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_830_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_829_wire_constant, tmp_var);
      EQ_u8_u1_830_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_834_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_833_wire_constant, tmp_var);
      EQ_u8_u1_834_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_838_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_837_wire_constant, tmp_var);
      EQ_u8_u1_838_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_842_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_841_wire_constant, tmp_var);
      EQ_u8_u1_842_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_846_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_845_wire_constant, tmp_var);
      EQ_u8_u1_846_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_850_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_849_wire_constant, tmp_var);
      EQ_u8_u1_850_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_854_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_853_wire_constant, tmp_var);
      EQ_u8_u1_854_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_858_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_857_wire_constant, tmp_var);
      EQ_u8_u1_858_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_862_inst
    process(op_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(op_560, konst_861_wire_constant, tmp_var);
      EQ_u8_u1_862_wire <= tmp_var; --
    end process;
    -- shared load operator group (0) : LOAD_next_pc1_795_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_next_pc1_795_load_0_req_0;
      LOAD_next_pc1_795_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_next_pc1_795_load_0_req_1;
      LOAD_next_pc1_795_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_next_pc1_795_word_address_0;
      LOAD_next_pc1_795_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(0 downto 0),
          mtag => memory_space_1_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(7 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : STORE_next_pc1_675_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_next_pc1_675_store_0_req_0;
      STORE_next_pc1_675_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_next_pc1_675_store_0_req_1;
      STORE_next_pc1_675_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= halt1_577(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_next_pc1_675_word_address_0;
      data_in <= STORE_next_pc1_675_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(0 downto 0),
          mdata => memory_space_1_sr_data(7 downto 0),
          mtag => memory_space_1_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared call operator group (0) : call_stmt_667_call call_stmt_672_call 
    accessreg_call_group_0: Block -- 
      signal data_in: std_logic_vector(81 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_667_call_req_0;
      reqL_unguarded(0) <= call_stmt_672_call_req_0;
      call_stmt_667_call_ack_0 <= ackL_unguarded(1);
      call_stmt_672_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_667_call_req_1;
      reqR_unguarded(0) <= call_stmt_672_call_req_1;
      call_stmt_667_call_ack_1 <= ackR_unguarded(1);
      call_stmt_672_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessreg_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessreg_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessreg_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessreg_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessreg_call_group_0_gI: SplitGuardInterface generic map(name => "accessreg_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_663_wire_constant & rs1_564 & konst_665_wire_constant & konst_668_wire_constant & rs2_568 & konst_670_wire_constant;
      rs1_data_667 <= data_out(63 downto 32);
      rs2_data_672 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 82,
        owidth => 41,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessreg_call_reqs(0),
          ackR => accessreg_call_acks(0),
          dataR => accessreg_call_data(40 downto 0),
          tagR => accessreg_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessreg_return_acks(0), -- cross-over
          ackL => accessreg_return_reqs(0), -- cross-over
          dataL => accessreg_return_data(31 downto 0),
          tagL => accessreg_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_676_call 
    halt_call_group_1: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_676_call_req_0;
      call_stmt_676_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_676_call_req_1;
      call_stmt_676_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= halt1_577(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      halt_call_group_1_gI: SplitGuardInterface generic map(name => "halt_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= pc_buffer;
      STORE_next_pc1_675_wire <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 8,
        owidth => 8,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => halt_call_reqs(0),
          ackR => halt_call_acks(0),
          dataR => halt_call_data(7 downto 0),
          tagR => halt_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => halt_return_acks(0), -- cross-over
          ackL => halt_return_reqs(0), -- cross-over
          dataL => halt_return_data(7 downto 0),
          tagL => halt_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_682_call 
    sbir_call_group_2: Block -- 
      signal data_in: std_logic_vector(23 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_682_call_req_0;
      call_stmt_682_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_682_call_req_1;
      call_stmt_682_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= sbir1_582(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sbir_call_group_2_gI: SplitGuardInterface generic map(name => "sbir_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rs1_564 & rd_572 & pc_buffer;
      next_pc2_682 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 24,
        owidth => 24,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => sbir_call_reqs(0),
          ackR => sbir_call_acks(0),
          dataR => sbir_call_data(23 downto 0),
          tagR => sbir_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => sbir_return_acks(0), -- cross-over
          ackL => sbir_return_reqs(0), -- cross-over
          dataL => sbir_return_data(7 downto 0),
          tagL => sbir_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_688_call 
    load_call_group_3: Block -- 
      signal data_in: std_logic_vector(47 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_688_call_req_0;
      call_stmt_688_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_688_call_req_1;
      call_stmt_688_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= load1_587(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      load_call_group_3_gI: SplitGuardInterface generic map(name => "load_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rs1_data_667 & rd_572 & pc_buffer;
      next_pc3_688 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 48,
        owidth => 48,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => load_call_reqs(0),
          ackR => load_call_acks(0),
          dataR => load_call_data(47 downto 0),
          tagR => load_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => load_return_acks(0), -- cross-over
          ackL => load_return_reqs(0), -- cross-over
          dataL => load_return_data(7 downto 0),
          tagL => load_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- shared call operator group (4) : call_stmt_694_call 
    store_call_group_4: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_694_call_req_0;
      call_stmt_694_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_694_call_req_1;
      call_stmt_694_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= store1_592(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      store_call_group_4_gI: SplitGuardInterface generic map(name => "store_call_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rs1_data_667 & rs2_data_672 & pc_buffer;
      next_pc4_694 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 72,
        owidth => 72,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => store_call_reqs(0),
          ackR => store_call_acks(0),
          dataR => store_call_data(71 downto 0),
          tagR => store_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => store_return_acks(0), -- cross-over
          ackL => store_return_reqs(0), -- cross-over
          dataL => store_return_data(7 downto 0),
          tagL => store_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    -- shared call operator group (5) : call_stmt_701_call 
    and_i_call_group_5: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_701_call_req_0;
      call_stmt_701_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_701_call_req_1;
      call_stmt_701_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= and1_597(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      and_i_call_group_5_gI: SplitGuardInterface generic map(name => "and_i_call_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rs1_data_667 & rs2_data_672 & rd_572 & pc_buffer;
      next_pc5_701 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 80,
        owidth => 80,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => and_i_call_reqs(0),
          ackR => and_i_call_acks(0),
          dataR => and_i_call_data(79 downto 0),
          tagR => and_i_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => and_i_return_acks(0), -- cross-over
          ackL => and_i_return_reqs(0), -- cross-over
          dataL => and_i_return_data(7 downto 0),
          tagL => and_i_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 5
    -- shared call operator group (6) : call_stmt_708_call 
    or_i_call_group_6: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_708_call_req_0;
      call_stmt_708_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_708_call_req_1;
      call_stmt_708_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= or1_602(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      or_i_call_group_6_gI: SplitGuardInterface generic map(name => "or_i_call_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rs1_data_667 & rs2_data_672 & rd_572 & pc_buffer;
      next_pc6_708 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 80,
        owidth => 80,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => or_i_call_reqs(0),
          ackR => or_i_call_acks(0),
          dataR => or_i_call_data(79 downto 0),
          tagR => or_i_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => or_i_return_acks(0), -- cross-over
          ackL => or_i_return_reqs(0), -- cross-over
          dataL => or_i_return_data(7 downto 0),
          tagL => or_i_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 6
    -- shared call operator group (7) : call_stmt_715_call 
    xnor_i_call_group_7: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_715_call_req_0;
      call_stmt_715_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_715_call_req_1;
      call_stmt_715_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= xnor1_607(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      xnor_i_call_group_7_gI: SplitGuardInterface generic map(name => "xnor_i_call_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rs1_data_667 & rs2_data_672 & rd_572 & pc_buffer;
      next_pc7_715 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 80,
        owidth => 80,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => xnor_i_call_reqs(0),
          ackR => xnor_i_call_acks(0),
          dataR => xnor_i_call_data(79 downto 0),
          tagR => xnor_i_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => xnor_i_return_acks(0), -- cross-over
          ackL => xnor_i_return_reqs(0), -- cross-over
          dataL => xnor_i_return_data(7 downto 0),
          tagL => xnor_i_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 7
    -- shared call operator group (8) : call_stmt_722_call 
    xor_i_call_group_8: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_722_call_req_0;
      call_stmt_722_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_722_call_req_1;
      call_stmt_722_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= xor1_612(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      xor_i_call_group_8_gI: SplitGuardInterface generic map(name => "xor_i_call_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rs1_data_667 & rs2_data_672 & rd_572 & pc_buffer;
      next_pc8_722 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 80,
        owidth => 80,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => xor_i_call_reqs(0),
          ackR => xor_i_call_acks(0),
          dataR => xor_i_call_data(79 downto 0),
          tagR => xor_i_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => xor_i_return_acks(0), -- cross-over
          ackL => xor_i_return_reqs(0), -- cross-over
          dataL => xor_i_return_data(7 downto 0),
          tagL => xor_i_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 8
    -- shared call operator group (9) : call_stmt_729_call 
    add_call_group_9: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_729_call_req_0;
      call_stmt_729_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_729_call_req_1;
      call_stmt_729_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= add1_617(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      add_call_group_9_gI: SplitGuardInterface generic map(name => "add_call_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rs1_data_667 & rs2_data_672 & rd_572 & pc_buffer;
      next_pc9_729 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 80,
        owidth => 80,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => add_call_reqs(0),
          ackR => add_call_acks(0),
          dataR => add_call_data(79 downto 0),
          tagR => add_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => add_return_acks(0), -- cross-over
          ackL => add_return_reqs(0), -- cross-over
          dataL => add_return_data(7 downto 0),
          tagL => add_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 9
    -- shared call operator group (10) : call_stmt_736_call 
    sub_call_group_10: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_736_call_req_0;
      call_stmt_736_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_736_call_req_1;
      call_stmt_736_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= sub1_622(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sub_call_group_10_gI: SplitGuardInterface generic map(name => "sub_call_group_10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rs1_data_667 & rs2_data_672 & rd_572 & pc_buffer;
      next_pc10_736 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 80,
        owidth => 80,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => sub_call_reqs(0),
          ackR => sub_call_acks(0),
          dataR => sub_call_data(79 downto 0),
          tagR => sub_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => sub_return_acks(0), -- cross-over
          ackL => sub_return_reqs(0), -- cross-over
          dataL => sub_return_data(7 downto 0),
          tagL => sub_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 10
    -- shared call operator group (11) : call_stmt_743_call 
    sll_i_call_group_11: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_743_call_req_0;
      call_stmt_743_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_743_call_req_1;
      call_stmt_743_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= sll1_627(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sll_i_call_group_11_gI: SplitGuardInterface generic map(name => "sll_i_call_group_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rs1_data_667 & rs2_data_672 & rd_572 & pc_buffer;
      next_pc11_743 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 80,
        owidth => 80,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => sll_i_call_reqs(0),
          ackR => sll_i_call_acks(0),
          dataR => sll_i_call_data(79 downto 0),
          tagR => sll_i_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => sll_i_return_acks(0), -- cross-over
          ackL => sll_i_return_reqs(0), -- cross-over
          dataL => sll_i_return_data(7 downto 0),
          tagL => sll_i_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 11
    -- shared call operator group (12) : call_stmt_750_call 
    srl_i_call_group_12: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_750_call_req_0;
      call_stmt_750_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_750_call_req_1;
      call_stmt_750_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= srl1_632(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      srl_i_call_group_12_gI: SplitGuardInterface generic map(name => "srl_i_call_group_12_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rs1_data_667 & rs2_data_672 & rd_572 & pc_buffer;
      next_pc12_750 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 80,
        owidth => 80,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => srl_i_call_reqs(0),
          ackR => srl_i_call_acks(0),
          dataR => srl_i_call_data(79 downto 0),
          tagR => srl_i_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => srl_i_return_acks(0), -- cross-over
          ackL => srl_i_return_reqs(0), -- cross-over
          dataL => srl_i_return_data(7 downto 0),
          tagL => srl_i_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 12
    -- shared call operator group (13) : call_stmt_757_call 
    sra_i_call_group_13: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_757_call_req_0;
      call_stmt_757_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_757_call_req_1;
      call_stmt_757_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= sra1_637(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sra_i_call_group_13_gI: SplitGuardInterface generic map(name => "sra_i_call_group_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rs1_data_667 & rs2_data_672 & rd_572 & pc_buffer;
      next_pc13_757 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 80,
        owidth => 80,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => sra_i_call_reqs(0),
          ackR => sra_i_call_acks(0),
          dataR => sra_i_call_data(79 downto 0),
          tagR => sra_i_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => sra_i_return_acks(0), -- cross-over
          ackL => sra_i_return_reqs(0), -- cross-over
          dataL => sra_i_return_data(7 downto 0),
          tagL => sra_i_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 13
    -- shared call operator group (14) : call_stmt_764_call 
    bz_call_group_14: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_764_call_req_0;
      call_stmt_764_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_764_call_req_1;
      call_stmt_764_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= bz1_642(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      bz_call_group_14_gI: SplitGuardInterface generic map(name => "bz_call_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rs1_data_667 & rs2_data_672 & rd_572 & pc_buffer;
      next_pc14_764 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 80,
        owidth => 80,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => bz_call_reqs(0),
          ackR => bz_call_acks(0),
          dataR => bz_call_data(79 downto 0),
          tagR => bz_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => bz_return_acks(0), -- cross-over
          ackL => bz_return_reqs(0), -- cross-over
          dataL => bz_return_data(7 downto 0),
          tagL => bz_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 14
    -- shared call operator group (15) : call_stmt_771_call 
    bn_call_group_15: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_771_call_req_0;
      call_stmt_771_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_771_call_req_1;
      call_stmt_771_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= bn1_647(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      bn_call_group_15_gI: SplitGuardInterface generic map(name => "bn_call_group_15_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rs1_data_667 & rs2_data_672 & rd_572 & pc_buffer;
      next_pc15_771 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 80,
        owidth => 80,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => bn_call_reqs(0),
          ackR => bn_call_acks(0),
          dataR => bn_call_data(79 downto 0),
          tagR => bn_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => bn_return_acks(0), -- cross-over
          ackL => bn_return_reqs(0), -- cross-over
          dataL => bn_return_data(7 downto 0),
          tagL => bn_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 15
    -- shared call operator group (16) : call_stmt_778_call 
    call_call_group_16: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_778_call_req_0;
      call_stmt_778_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_778_call_req_1;
      call_stmt_778_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= call1_652(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      call_call_group_16_gI: SplitGuardInterface generic map(name => "call_call_group_16_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rs1_data_667 & rs2_data_672 & rd_572 & pc_buffer;
      next_pc16_778 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 80,
        owidth => 80,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => call_call_reqs(0),
          ackR => call_call_acks(0),
          dataR => call_call_data(79 downto 0),
          tagR => call_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => call_return_acks(0), -- cross-over
          ackL => call_return_reqs(0), -- cross-over
          dataL => call_return_data(7 downto 0),
          tagL => call_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 16
    -- shared call operator group (17) : call_stmt_783_call 
    jmp_call_group_17: Block -- 
      signal data_in: std_logic_vector(39 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_783_call_req_0;
      call_stmt_783_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_783_call_req_1;
      call_stmt_783_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= jmp1_657(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      jmp_call_group_17_gI: SplitGuardInterface generic map(name => "jmp_call_group_17_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rs1_data_667 & pc_buffer;
      next_pc17_783 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 40,
        owidth => 40,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => jmp_call_reqs(0),
          ackR => jmp_call_acks(0),
          dataR => jmp_call_data(39 downto 0),
          tagR => jmp_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => jmp_return_acks(0), -- cross-over
          ackL => jmp_return_reqs(0), -- cross-over
          dataL => jmp_return_data(7 downto 0),
          tagL => jmp_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 17
    -- shared call operator group (18) : call_stmt_790_call 
    cmp_call_group_18: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_790_call_req_0;
      call_stmt_790_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_790_call_req_1;
      call_stmt_790_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= cmp1_662(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      cmp_call_group_18_gI: SplitGuardInterface generic map(name => "cmp_call_group_18_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rs1_data_667 & rs2_data_672 & rd_572 & pc_buffer;
      next_pc18_790 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 80,
        owidth => 80,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => cmp_call_reqs(0),
          ackR => cmp_call_acks(0),
          dataR => cmp_call_data(79 downto 0),
          tagR => cmp_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => cmp_return_acks(0), -- cross-over
          ackL => cmp_return_reqs(0), -- cross-over
          dataL => cmp_return_data(7 downto 0),
          tagL => cmp_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 18
    -- 
  end Block; -- data_path
  -- 
end try_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity try1 is -- 
  generic (tag_length : integer); 
  port ( -- 
    write_mem_pipe_read_req : out  std_logic_vector(0 downto 0);
    write_mem_pipe_read_ack : in   std_logic_vector(0 downto 0);
    write_mem_pipe_read_data : in   std_logic_vector(7 downto 0);
    LEDS_pipe_write_req : out  std_logic_vector(0 downto 0);
    LEDS_pipe_write_ack : in   std_logic_vector(0 downto 0);
    LEDS_pipe_write_data : out  std_logic_vector(15 downto 0);
    reg_output_pipe_write_req : out  std_logic_vector(0 downto 0);
    reg_output_pipe_write_ack : in   std_logic_vector(0 downto 0);
    reg_output_pipe_write_data : out  std_logic_vector(7 downto 0);
    init_mem_call_reqs : out  std_logic_vector(0 downto 0);
    init_mem_call_acks : in   std_logic_vector(0 downto 0);
    init_mem_call_tag  :  out  std_logic_vector(0 downto 0);
    init_mem_return_reqs : out  std_logic_vector(0 downto 0);
    init_mem_return_acks : in   std_logic_vector(0 downto 0);
    init_mem_return_tag :  in   std_logic_vector(0 downto 0);
    init_reg_call_reqs : out  std_logic_vector(0 downto 0);
    init_reg_call_acks : in   std_logic_vector(0 downto 0);
    init_reg_call_tag  :  out  std_logic_vector(0 downto 0);
    init_reg_return_reqs : out  std_logic_vector(0 downto 0);
    init_reg_return_acks : in   std_logic_vector(0 downto 0);
    init_reg_return_tag :  in   std_logic_vector(0 downto 0);
    try_call_reqs : out  std_logic_vector(0 downto 0);
    try_call_acks : in   std_logic_vector(0 downto 0);
    try_call_data : out  std_logic_vector(39 downto 0);
    try_call_tag  :  out  std_logic_vector(0 downto 0);
    try_return_reqs : out  std_logic_vector(0 downto 0);
    try_return_acks : in   std_logic_vector(0 downto 0);
    try_return_data : in   std_logic_vector(7 downto 0);
    try_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity try1;
architecture try1_arch of try1 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal try1_CP_2356_start: Boolean;
  signal try1_CP_2356_symbol: Boolean;
  -- volatile/operator module components. 
  component init_mem is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component init_reg is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component try is -- 
    generic (tag_length : integer); 
    port ( -- 
      pc : in  std_logic_vector(7 downto 0);
      inst : in  std_logic_vector(31 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      cmp_call_reqs : out  std_logic_vector(0 downto 0);
      cmp_call_acks : in   std_logic_vector(0 downto 0);
      cmp_call_data : out  std_logic_vector(79 downto 0);
      cmp_call_tag  :  out  std_logic_vector(0 downto 0);
      cmp_return_reqs : out  std_logic_vector(0 downto 0);
      cmp_return_acks : in   std_logic_vector(0 downto 0);
      cmp_return_data : in   std_logic_vector(7 downto 0);
      cmp_return_tag :  in   std_logic_vector(0 downto 0);
      sub_call_reqs : out  std_logic_vector(0 downto 0);
      sub_call_acks : in   std_logic_vector(0 downto 0);
      sub_call_data : out  std_logic_vector(79 downto 0);
      sub_call_tag  :  out  std_logic_vector(0 downto 0);
      sub_return_reqs : out  std_logic_vector(0 downto 0);
      sub_return_acks : in   std_logic_vector(0 downto 0);
      sub_return_data : in   std_logic_vector(7 downto 0);
      sub_return_tag :  in   std_logic_vector(0 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      bn_call_reqs : out  std_logic_vector(0 downto 0);
      bn_call_acks : in   std_logic_vector(0 downto 0);
      bn_call_data : out  std_logic_vector(79 downto 0);
      bn_call_tag  :  out  std_logic_vector(0 downto 0);
      bn_return_reqs : out  std_logic_vector(0 downto 0);
      bn_return_acks : in   std_logic_vector(0 downto 0);
      bn_return_data : in   std_logic_vector(7 downto 0);
      bn_return_tag :  in   std_logic_vector(0 downto 0);
      halt_call_reqs : out  std_logic_vector(0 downto 0);
      halt_call_acks : in   std_logic_vector(0 downto 0);
      halt_call_data : out  std_logic_vector(7 downto 0);
      halt_call_tag  :  out  std_logic_vector(0 downto 0);
      halt_return_reqs : out  std_logic_vector(0 downto 0);
      halt_return_acks : in   std_logic_vector(0 downto 0);
      halt_return_data : in   std_logic_vector(7 downto 0);
      halt_return_tag :  in   std_logic_vector(0 downto 0);
      add_call_reqs : out  std_logic_vector(0 downto 0);
      add_call_acks : in   std_logic_vector(0 downto 0);
      add_call_data : out  std_logic_vector(79 downto 0);
      add_call_tag  :  out  std_logic_vector(0 downto 0);
      add_return_reqs : out  std_logic_vector(0 downto 0);
      add_return_acks : in   std_logic_vector(0 downto 0);
      add_return_data : in   std_logic_vector(7 downto 0);
      add_return_tag :  in   std_logic_vector(0 downto 0);
      sll_i_call_reqs : out  std_logic_vector(0 downto 0);
      sll_i_call_acks : in   std_logic_vector(0 downto 0);
      sll_i_call_data : out  std_logic_vector(79 downto 0);
      sll_i_call_tag  :  out  std_logic_vector(0 downto 0);
      sll_i_return_reqs : out  std_logic_vector(0 downto 0);
      sll_i_return_acks : in   std_logic_vector(0 downto 0);
      sll_i_return_data : in   std_logic_vector(7 downto 0);
      sll_i_return_tag :  in   std_logic_vector(0 downto 0);
      and_i_call_reqs : out  std_logic_vector(0 downto 0);
      and_i_call_acks : in   std_logic_vector(0 downto 0);
      and_i_call_data : out  std_logic_vector(79 downto 0);
      and_i_call_tag  :  out  std_logic_vector(0 downto 0);
      and_i_return_reqs : out  std_logic_vector(0 downto 0);
      and_i_return_acks : in   std_logic_vector(0 downto 0);
      and_i_return_data : in   std_logic_vector(7 downto 0);
      and_i_return_tag :  in   std_logic_vector(0 downto 0);
      call_call_reqs : out  std_logic_vector(0 downto 0);
      call_call_acks : in   std_logic_vector(0 downto 0);
      call_call_data : out  std_logic_vector(79 downto 0);
      call_call_tag  :  out  std_logic_vector(0 downto 0);
      call_return_reqs : out  std_logic_vector(0 downto 0);
      call_return_acks : in   std_logic_vector(0 downto 0);
      call_return_data : in   std_logic_vector(7 downto 0);
      call_return_tag :  in   std_logic_vector(0 downto 0);
      bz_call_reqs : out  std_logic_vector(0 downto 0);
      bz_call_acks : in   std_logic_vector(0 downto 0);
      bz_call_data : out  std_logic_vector(79 downto 0);
      bz_call_tag  :  out  std_logic_vector(0 downto 0);
      bz_return_reqs : out  std_logic_vector(0 downto 0);
      bz_return_acks : in   std_logic_vector(0 downto 0);
      bz_return_data : in   std_logic_vector(7 downto 0);
      bz_return_tag :  in   std_logic_vector(0 downto 0);
      xnor_i_call_reqs : out  std_logic_vector(0 downto 0);
      xnor_i_call_acks : in   std_logic_vector(0 downto 0);
      xnor_i_call_data : out  std_logic_vector(79 downto 0);
      xnor_i_call_tag  :  out  std_logic_vector(0 downto 0);
      xnor_i_return_reqs : out  std_logic_vector(0 downto 0);
      xnor_i_return_acks : in   std_logic_vector(0 downto 0);
      xnor_i_return_data : in   std_logic_vector(7 downto 0);
      xnor_i_return_tag :  in   std_logic_vector(0 downto 0);
      sra_i_call_reqs : out  std_logic_vector(0 downto 0);
      sra_i_call_acks : in   std_logic_vector(0 downto 0);
      sra_i_call_data : out  std_logic_vector(79 downto 0);
      sra_i_call_tag  :  out  std_logic_vector(0 downto 0);
      sra_i_return_reqs : out  std_logic_vector(0 downto 0);
      sra_i_return_acks : in   std_logic_vector(0 downto 0);
      sra_i_return_data : in   std_logic_vector(7 downto 0);
      sra_i_return_tag :  in   std_logic_vector(0 downto 0);
      sbir_call_reqs : out  std_logic_vector(0 downto 0);
      sbir_call_acks : in   std_logic_vector(0 downto 0);
      sbir_call_data : out  std_logic_vector(23 downto 0);
      sbir_call_tag  :  out  std_logic_vector(0 downto 0);
      sbir_return_reqs : out  std_logic_vector(0 downto 0);
      sbir_return_acks : in   std_logic_vector(0 downto 0);
      sbir_return_data : in   std_logic_vector(7 downto 0);
      sbir_return_tag :  in   std_logic_vector(0 downto 0);
      or_i_call_reqs : out  std_logic_vector(0 downto 0);
      or_i_call_acks : in   std_logic_vector(0 downto 0);
      or_i_call_data : out  std_logic_vector(79 downto 0);
      or_i_call_tag  :  out  std_logic_vector(0 downto 0);
      or_i_return_reqs : out  std_logic_vector(0 downto 0);
      or_i_return_acks : in   std_logic_vector(0 downto 0);
      or_i_return_data : in   std_logic_vector(7 downto 0);
      or_i_return_tag :  in   std_logic_vector(0 downto 0);
      load_call_reqs : out  std_logic_vector(0 downto 0);
      load_call_acks : in   std_logic_vector(0 downto 0);
      load_call_data : out  std_logic_vector(47 downto 0);
      load_call_tag  :  out  std_logic_vector(0 downto 0);
      load_return_reqs : out  std_logic_vector(0 downto 0);
      load_return_acks : in   std_logic_vector(0 downto 0);
      load_return_data : in   std_logic_vector(7 downto 0);
      load_return_tag :  in   std_logic_vector(0 downto 0);
      jmp_call_reqs : out  std_logic_vector(0 downto 0);
      jmp_call_acks : in   std_logic_vector(0 downto 0);
      jmp_call_data : out  std_logic_vector(39 downto 0);
      jmp_call_tag  :  out  std_logic_vector(0 downto 0);
      jmp_return_reqs : out  std_logic_vector(0 downto 0);
      jmp_return_acks : in   std_logic_vector(0 downto 0);
      jmp_return_data : in   std_logic_vector(7 downto 0);
      jmp_return_tag :  in   std_logic_vector(0 downto 0);
      store_call_reqs : out  std_logic_vector(0 downto 0);
      store_call_acks : in   std_logic_vector(0 downto 0);
      store_call_data : out  std_logic_vector(71 downto 0);
      store_call_tag  :  out  std_logic_vector(0 downto 0);
      store_return_reqs : out  std_logic_vector(0 downto 0);
      store_return_acks : in   std_logic_vector(0 downto 0);
      store_return_data : in   std_logic_vector(7 downto 0);
      store_return_tag :  in   std_logic_vector(0 downto 0);
      srl_i_call_reqs : out  std_logic_vector(0 downto 0);
      srl_i_call_acks : in   std_logic_vector(0 downto 0);
      srl_i_call_data : out  std_logic_vector(79 downto 0);
      srl_i_call_tag  :  out  std_logic_vector(0 downto 0);
      srl_i_return_reqs : out  std_logic_vector(0 downto 0);
      srl_i_return_acks : in   std_logic_vector(0 downto 0);
      srl_i_return_data : in   std_logic_vector(7 downto 0);
      srl_i_return_tag :  in   std_logic_vector(0 downto 0);
      xor_i_call_reqs : out  std_logic_vector(0 downto 0);
      xor_i_call_acks : in   std_logic_vector(0 downto 0);
      xor_i_call_data : out  std_logic_vector(79 downto 0);
      xor_i_call_tag  :  out  std_logic_vector(0 downto 0);
      xor_i_return_reqs : out  std_logic_vector(0 downto 0);
      xor_i_return_acks : in   std_logic_vector(0 downto 0);
      xor_i_return_data : in   std_logic_vector(7 downto 0);
      xor_i_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_890_call_req_0 : boolean;
  signal call_stmt_890_call_ack_0 : boolean;
  signal call_stmt_890_call_req_1 : boolean;
  signal call_stmt_890_call_ack_1 : boolean;
  signal call_stmt_891_call_req_0 : boolean;
  signal call_stmt_891_call_ack_0 : boolean;
  signal call_stmt_891_call_req_1 : boolean;
  signal call_stmt_891_call_ack_1 : boolean;
  signal RPIPE_write_mem_901_inst_req_0 : boolean;
  signal RPIPE_write_mem_901_inst_ack_0 : boolean;
  signal RPIPE_write_mem_901_inst_req_1 : boolean;
  signal RPIPE_write_mem_901_inst_ack_1 : boolean;
  signal RPIPE_write_mem_904_inst_req_0 : boolean;
  signal RPIPE_write_mem_904_inst_ack_0 : boolean;
  signal RPIPE_write_mem_904_inst_req_1 : boolean;
  signal RPIPE_write_mem_904_inst_ack_1 : boolean;
  signal RPIPE_write_mem_907_inst_req_0 : boolean;
  signal RPIPE_write_mem_907_inst_ack_0 : boolean;
  signal RPIPE_write_mem_907_inst_req_1 : boolean;
  signal RPIPE_write_mem_907_inst_ack_1 : boolean;
  signal RPIPE_write_mem_910_inst_req_0 : boolean;
  signal RPIPE_write_mem_910_inst_ack_0 : boolean;
  signal RPIPE_write_mem_910_inst_req_1 : boolean;
  signal RPIPE_write_mem_910_inst_ack_1 : boolean;
  signal CONCAT_u16_u32_919_inst_req_0 : boolean;
  signal CONCAT_u16_u32_919_inst_ack_0 : boolean;
  signal CONCAT_u16_u32_919_inst_req_1 : boolean;
  signal CONCAT_u16_u32_919_inst_ack_1 : boolean;
  signal call_stmt_924_call_req_0 : boolean;
  signal call_stmt_924_call_ack_0 : boolean;
  signal call_stmt_924_call_req_1 : boolean;
  signal call_stmt_924_call_ack_1 : boolean;
  signal WPIPE_reg_output_925_inst_req_0 : boolean;
  signal WPIPE_reg_output_925_inst_ack_0 : boolean;
  signal WPIPE_reg_output_925_inst_req_1 : boolean;
  signal WPIPE_reg_output_925_inst_ack_1 : boolean;
  signal CONCAT_u8_u16_931_inst_req_0 : boolean;
  signal CONCAT_u8_u16_931_inst_ack_0 : boolean;
  signal CONCAT_u8_u16_931_inst_req_1 : boolean;
  signal CONCAT_u8_u16_931_inst_ack_1 : boolean;
  signal WPIPE_LEDS_928_inst_req_0 : boolean;
  signal WPIPE_LEDS_928_inst_ack_0 : boolean;
  signal WPIPE_LEDS_928_inst_req_1 : boolean;
  signal WPIPE_LEDS_928_inst_ack_1 : boolean;
  signal phi_stmt_894_req_0 : boolean;
  signal next_pc_924_898_buf_req_0 : boolean;
  signal next_pc_924_898_buf_ack_0 : boolean;
  signal next_pc_924_898_buf_req_1 : boolean;
  signal next_pc_924_898_buf_ack_1 : boolean;
  signal phi_stmt_894_req_1 : boolean;
  signal phi_stmt_894_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "try1_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  try1_CP_2356_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "try1_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= try1_CP_2356_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= try1_CP_2356_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= try1_CP_2356_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  try1_CP_2356: Block -- control-path 
    signal try1_CP_2356_elements: BooleanArray(33 downto 0);
    -- 
  begin -- 
    try1_CP_2356_elements(0) <= try1_CP_2356_start;
    try1_CP_2356_symbol <= try1_CP_2356_elements(6);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_890_to_call_stmt_891/$entry
      -- CP-element group 0: 	 call_stmt_890_to_call_stmt_891/call_stmt_890_sample_start_
      -- CP-element group 0: 	 call_stmt_890_to_call_stmt_891/call_stmt_890_update_start_
      -- CP-element group 0: 	 call_stmt_890_to_call_stmt_891/call_stmt_890_Sample/$entry
      -- CP-element group 0: 	 call_stmt_890_to_call_stmt_891/call_stmt_890_Sample/crr
      -- CP-element group 0: 	 call_stmt_890_to_call_stmt_891/call_stmt_890_Update/$entry
      -- CP-element group 0: 	 call_stmt_890_to_call_stmt_891/call_stmt_890_Update/ccr
      -- CP-element group 0: 	 call_stmt_890_to_call_stmt_891/call_stmt_891_sample_start_
      -- CP-element group 0: 	 call_stmt_890_to_call_stmt_891/call_stmt_891_update_start_
      -- CP-element group 0: 	 call_stmt_890_to_call_stmt_891/call_stmt_891_Sample/$entry
      -- CP-element group 0: 	 call_stmt_890_to_call_stmt_891/call_stmt_891_Sample/crr
      -- CP-element group 0: 	 call_stmt_890_to_call_stmt_891/call_stmt_891_Update/$entry
      -- CP-element group 0: 	 call_stmt_890_to_call_stmt_891/call_stmt_891_Update/ccr
      -- 
    crr_2369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(0), ack => call_stmt_890_call_req_0); -- 
    ccr_2374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(0), ack => call_stmt_890_call_req_1); -- 
    crr_2383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(0), ack => call_stmt_891_call_req_0); -- 
    ccr_2388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(0), ack => call_stmt_891_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_890_to_call_stmt_891/call_stmt_890_sample_completed_
      -- CP-element group 1: 	 call_stmt_890_to_call_stmt_891/call_stmt_890_Sample/$exit
      -- CP-element group 1: 	 call_stmt_890_to_call_stmt_891/call_stmt_890_Sample/cra
      -- 
    cra_2370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_890_call_ack_0, ack => try1_CP_2356_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 call_stmt_890_to_call_stmt_891/call_stmt_890_update_completed_
      -- CP-element group 2: 	 call_stmt_890_to_call_stmt_891/call_stmt_890_Update/$exit
      -- CP-element group 2: 	 call_stmt_890_to_call_stmt_891/call_stmt_890_Update/cca
      -- 
    cca_2375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_890_call_ack_1, ack => try1_CP_2356_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_890_to_call_stmt_891/call_stmt_891_sample_completed_
      -- CP-element group 3: 	 call_stmt_890_to_call_stmt_891/call_stmt_891_Sample/$exit
      -- CP-element group 3: 	 call_stmt_890_to_call_stmt_891/call_stmt_891_Sample/cra
      -- 
    cra_2384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_891_call_ack_0, ack => try1_CP_2356_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 call_stmt_890_to_call_stmt_891/call_stmt_891_update_completed_
      -- CP-element group 4: 	 call_stmt_890_to_call_stmt_891/call_stmt_891_Update/$exit
      -- CP-element group 4: 	 call_stmt_890_to_call_stmt_891/call_stmt_891_Update/cca
      -- 
    cca_2389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_891_call_ack_1, ack => try1_CP_2356_elements(4)); -- 
    -- CP-element group 5:  branch  join  transition  place  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	28 
    -- CP-element group 5:  members (8) 
      -- CP-element group 5: 	 call_stmt_890_to_call_stmt_891/$exit
      -- CP-element group 5: 	 branch_block_stmt_892/$entry
      -- CP-element group 5: 	 branch_block_stmt_892/branch_block_stmt_892__entry__
      -- CP-element group 5: 	 branch_block_stmt_892/merge_stmt_893__entry__
      -- CP-element group 5: 	 branch_block_stmt_892/merge_stmt_893_dead_link/$entry
      -- CP-element group 5: 	 branch_block_stmt_892/merge_stmt_893__entry___PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_892/merge_stmt_893__entry___PhiReq/phi_stmt_894/$entry
      -- CP-element group 5: 	 branch_block_stmt_892/merge_stmt_893__entry___PhiReq/phi_stmt_894/phi_stmt_894_sources/$entry
      -- 
    try1_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 23) := "try1_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_2356_elements(2) & try1_CP_2356_elements(4);
      gj_try1_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_2356_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  transition  place  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 $exit
      -- CP-element group 6: 	 branch_block_stmt_892/$exit
      -- CP-element group 6: 	 branch_block_stmt_892/branch_block_stmt_892__exit__
      -- 
    try1_CP_2356_elements(6) <= false; 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	33 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_901_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_901_update_start_
      -- CP-element group 7: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_901_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_901_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_901_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_901_Update/cr
      -- 
    ra_2411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_write_mem_901_inst_ack_0, ack => try1_CP_2356_elements(7)); -- 
    cr_2415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(7), ack => RPIPE_write_mem_901_inst_req_1); -- 
    -- CP-element group 8:  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	15 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_901_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_901_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_901_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_904_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_904_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_904_Sample/rr
      -- 
    ca_2416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_write_mem_901_inst_ack_1, ack => try1_CP_2356_elements(8)); -- 
    rr_2424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(8), ack => RPIPE_write_mem_904_inst_req_0); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_904_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_904_update_start_
      -- CP-element group 9: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_904_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_904_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_904_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_904_Update/cr
      -- 
    ra_2425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_write_mem_904_inst_ack_0, ack => try1_CP_2356_elements(9)); -- 
    cr_2429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(9), ack => RPIPE_write_mem_904_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_904_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_904_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_904_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_907_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_907_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_907_Sample/rr
      -- 
    ca_2430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_write_mem_904_inst_ack_1, ack => try1_CP_2356_elements(10)); -- 
    rr_2438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(10), ack => RPIPE_write_mem_907_inst_req_0); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_907_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_907_update_start_
      -- CP-element group 11: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_907_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_907_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_907_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_907_Update/cr
      -- 
    ra_2439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_write_mem_907_inst_ack_0, ack => try1_CP_2356_elements(11)); -- 
    cr_2443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(11), ack => RPIPE_write_mem_907_inst_req_1); -- 
    -- CP-element group 12:  fork  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_907_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_907_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_907_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_910_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_910_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_910_Sample/rr
      -- 
    ca_2444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_write_mem_907_inst_ack_1, ack => try1_CP_2356_elements(12)); -- 
    rr_2452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(12), ack => RPIPE_write_mem_910_inst_req_0); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_910_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_910_update_start_
      -- CP-element group 13: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_910_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_910_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_910_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_910_Update/cr
      -- 
    ra_2453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_write_mem_910_inst_ack_0, ack => try1_CP_2356_elements(13)); -- 
    cr_2457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(13), ack => RPIPE_write_mem_910_inst_req_1); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_910_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_910_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_910_Update/ca
      -- 
    ca_2458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_write_mem_910_inst_ack_1, ack => try1_CP_2356_elements(14)); -- 
    -- CP-element group 15:  join  transition  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: 	10 
    -- CP-element group 15: 	12 
    -- CP-element group 15: 	8 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u16_u32_919_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u16_u32_919_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u16_u32_919_Sample/rr
      -- 
    rr_2466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(15), ack => CONCAT_u16_u32_919_inst_req_0); -- 
    try1_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= try1_CP_2356_elements(14) & try1_CP_2356_elements(10) & try1_CP_2356_elements(12) & try1_CP_2356_elements(8);
      gj_try1_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_2356_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u16_u32_919_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u16_u32_919_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u16_u32_919_Sample/ra
      -- 
    ra_2467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_919_inst_ack_0, ack => try1_CP_2356_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	33 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u16_u32_919_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u16_u32_919_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u16_u32_919_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/call_stmt_924_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/call_stmt_924_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/call_stmt_924_Sample/crr
      -- 
    ca_2472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_919_inst_ack_1, ack => try1_CP_2356_elements(17)); -- 
    crr_2480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(17), ack => call_stmt_924_call_req_0); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/call_stmt_924_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/call_stmt_924_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/call_stmt_924_Sample/cra
      -- 
    cra_2481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_924_call_ack_0, ack => try1_CP_2356_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	33 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/call_stmt_924_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/call_stmt_924_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/call_stmt_924_Update/cca
      -- 
    cca_2486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_924_call_ack_1, ack => try1_CP_2356_elements(19)); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	22 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_reg_output_925_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_reg_output_925_update_start_
      -- CP-element group 20: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_reg_output_925_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_reg_output_925_Sample/ack
      -- CP-element group 20: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_reg_output_925_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_reg_output_925_Update/req
      -- 
    ack_2495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_reg_output_925_inst_ack_0, ack => try1_CP_2356_elements(20)); -- 
    req_2499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(20), ack => WPIPE_reg_output_925_inst_req_1); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	27 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_reg_output_925_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_reg_output_925_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_reg_output_925_Update/ack
      -- 
    ack_2500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_reg_output_925_inst_ack_1, ack => try1_CP_2356_elements(21)); -- 
    -- CP-element group 22:  transition  output  delay-element  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	20 
    -- CP-element group 22:  members (4) 
      -- CP-element group 22: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_reg_output_925_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_reg_output_925_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_reg_output_925_Sample/req
      -- CP-element group 22: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/synch_WPIPE_reg_output_925_sample_start__call_stmt_924_sample_completed_
      -- 
    req_2494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(22), ack => WPIPE_reg_output_925_inst_req_0); -- 
    -- Element group try1_CP_2356_elements(22) is a control-delay.
    cp_element_22_delay: control_delay_element  generic map(name => " 22_delay", delay_value => 1)  port map(req => try1_CP_2356_elements(19), ack => try1_CP_2356_elements(22), clk => clk, reset =>reset);
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	33 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u8_u16_931_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u8_u16_931_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u8_u16_931_Sample/ra
      -- 
    ra_2510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u8_u16_931_inst_ack_0, ack => try1_CP_2356_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	33 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u8_u16_931_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u8_u16_931_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u8_u16_931_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_LEDS_928_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_LEDS_928_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_LEDS_928_Sample/req
      -- 
    ca_2515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u8_u16_931_inst_ack_1, ack => try1_CP_2356_elements(24)); -- 
    req_2523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(24), ack => WPIPE_LEDS_928_inst_req_0); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_LEDS_928_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_LEDS_928_update_start_
      -- CP-element group 25: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_LEDS_928_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_LEDS_928_Sample/ack
      -- CP-element group 25: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_LEDS_928_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_LEDS_928_Update/req
      -- 
    ack_2524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LEDS_928_inst_ack_0, ack => try1_CP_2356_elements(25)); -- 
    req_2528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(25), ack => WPIPE_LEDS_928_inst_req_1); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_LEDS_928_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_LEDS_928_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/WPIPE_LEDS_928_Update/ack
      -- 
    ack_2529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LEDS_928_inst_ack_1, ack => try1_CP_2356_elements(26)); -- 
    -- CP-element group 27:  join  fork  transition  place  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: 	21 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: 	30 
    -- CP-element group 27:  members (11) 
      -- CP-element group 27: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932__exit__
      -- CP-element group 27: 	 branch_block_stmt_892/loopback
      -- CP-element group 27: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/$exit
      -- CP-element group 27: 	 branch_block_stmt_892/loopback_PhiReq/$entry
      -- CP-element group 27: 	 branch_block_stmt_892/loopback_PhiReq/phi_stmt_894/$entry
      -- CP-element group 27: 	 branch_block_stmt_892/loopback_PhiReq/phi_stmt_894/phi_stmt_894_sources/$entry
      -- CP-element group 27: 	 branch_block_stmt_892/loopback_PhiReq/phi_stmt_894/phi_stmt_894_sources/Interlock/$entry
      -- CP-element group 27: 	 branch_block_stmt_892/loopback_PhiReq/phi_stmt_894/phi_stmt_894_sources/Interlock/Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_892/loopback_PhiReq/phi_stmt_894/phi_stmt_894_sources/Interlock/Sample/req
      -- CP-element group 27: 	 branch_block_stmt_892/loopback_PhiReq/phi_stmt_894/phi_stmt_894_sources/Interlock/Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_892/loopback_PhiReq/phi_stmt_894/phi_stmt_894_sources/Interlock/Update/req
      -- 
    req_2560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(27), ack => next_pc_924_898_buf_req_0); -- 
    req_2565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(27), ack => next_pc_924_898_buf_req_1); -- 
    try1_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_2356_elements(26) & try1_CP_2356_elements(21);
      gj_try1_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_2356_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  transition  output  delay-element  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	5 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	32 
    -- CP-element group 28:  members (5) 
      -- CP-element group 28: 	 branch_block_stmt_892/merge_stmt_893__entry___PhiReq/$exit
      -- CP-element group 28: 	 branch_block_stmt_892/merge_stmt_893__entry___PhiReq/phi_stmt_894/$exit
      -- CP-element group 28: 	 branch_block_stmt_892/merge_stmt_893__entry___PhiReq/phi_stmt_894/phi_stmt_894_sources/$exit
      -- CP-element group 28: 	 branch_block_stmt_892/merge_stmt_893__entry___PhiReq/phi_stmt_894/phi_stmt_894_sources/type_cast_897_konst_delay_trans
      -- CP-element group 28: 	 branch_block_stmt_892/merge_stmt_893__entry___PhiReq/phi_stmt_894/phi_stmt_894_req
      -- 
    phi_stmt_894_req_2544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_894_req_2544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(28), ack => phi_stmt_894_req_0); -- 
    -- Element group try1_CP_2356_elements(28) is a control-delay.
    cp_element_28_delay: control_delay_element  generic map(name => " 28_delay", delay_value => 1)  port map(req => try1_CP_2356_elements(5), ack => try1_CP_2356_elements(28), clk => clk, reset =>reset);
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_892/loopback_PhiReq/phi_stmt_894/phi_stmt_894_sources/Interlock/Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_892/loopback_PhiReq/phi_stmt_894/phi_stmt_894_sources/Interlock/Sample/ack
      -- 
    ack_2561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pc_924_898_buf_ack_0, ack => try1_CP_2356_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_892/loopback_PhiReq/phi_stmt_894/phi_stmt_894_sources/Interlock/Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_892/loopback_PhiReq/phi_stmt_894/phi_stmt_894_sources/Interlock/Update/ack
      -- 
    ack_2566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pc_924_898_buf_ack_1, ack => try1_CP_2356_elements(30)); -- 
    -- CP-element group 31:  join  transition  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (5) 
      -- CP-element group 31: 	 branch_block_stmt_892/loopback_PhiReq/$exit
      -- CP-element group 31: 	 branch_block_stmt_892/loopback_PhiReq/phi_stmt_894/$exit
      -- CP-element group 31: 	 branch_block_stmt_892/loopback_PhiReq/phi_stmt_894/phi_stmt_894_sources/$exit
      -- CP-element group 31: 	 branch_block_stmt_892/loopback_PhiReq/phi_stmt_894/phi_stmt_894_sources/Interlock/$exit
      -- CP-element group 31: 	 branch_block_stmt_892/loopback_PhiReq/phi_stmt_894/phi_stmt_894_req
      -- 
    phi_stmt_894_req_2567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_894_req_2567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(31), ack => phi_stmt_894_req_1); -- 
    try1_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "try1_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= try1_CP_2356_elements(29) & try1_CP_2356_elements(30);
      gj_try1_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => try1_CP_2356_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  merge  transition  place  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: 	28 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_892/merge_stmt_893_PhiReqMerge
      -- CP-element group 32: 	 branch_block_stmt_892/merge_stmt_893_PhiAck/$entry
      -- 
    try1_CP_2356_elements(32) <= OrReduce(try1_CP_2356_elements(31) & try1_CP_2356_elements(28));
    -- CP-element group 33:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	23 
    -- CP-element group 33: 	24 
    -- CP-element group 33: 	19 
    -- CP-element group 33: 	17 
    -- CP-element group 33: 	7 
    -- CP-element group 33:  members (20) 
      -- CP-element group 33: 	 branch_block_stmt_892/merge_stmt_893__exit__
      -- CP-element group 33: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932__entry__
      -- CP-element group 33: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/$entry
      -- CP-element group 33: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_901_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_901_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/RPIPE_write_mem_901_Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u16_u32_919_update_start_
      -- CP-element group 33: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u16_u32_919_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u16_u32_919_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/call_stmt_924_update_start_
      -- CP-element group 33: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/call_stmt_924_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/call_stmt_924_Update/ccr
      -- CP-element group 33: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u8_u16_931_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u8_u16_931_update_start_
      -- CP-element group 33: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u8_u16_931_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u8_u16_931_Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u8_u16_931_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_892/assign_stmt_902_to_assign_stmt_932/CONCAT_u8_u16_931_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_892/merge_stmt_893_PhiAck/$exit
      -- CP-element group 33: 	 branch_block_stmt_892/merge_stmt_893_PhiAck/phi_stmt_894_ack
      -- 
    phi_stmt_894_ack_2572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_894_ack_0, ack => try1_CP_2356_elements(33)); -- 
    rr_2410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(33), ack => RPIPE_write_mem_901_inst_req_0); -- 
    cr_2471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(33), ack => CONCAT_u16_u32_919_inst_req_1); -- 
    ccr_2485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(33), ack => call_stmt_924_call_req_1); -- 
    rr_2509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(33), ack => CONCAT_u8_u16_931_inst_req_0); -- 
    cr_2514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => try1_CP_2356_elements(33), ack => CONCAT_u8_u16_931_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u8_u16_915_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_918_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_931_wire : std_logic_vector(15 downto 0);
    signal R_zero8_929_wire_constant : std_logic_vector(7 downto 0);
    signal inst1_902 : std_logic_vector(7 downto 0);
    signal inst2_905 : std_logic_vector(7 downto 0);
    signal inst3_908 : std_logic_vector(7 downto 0);
    signal inst4_911 : std_logic_vector(7 downto 0);
    signal inst_920 : std_logic_vector(31 downto 0);
    signal next_pc_924 : std_logic_vector(7 downto 0);
    signal next_pc_924_898_buffered : std_logic_vector(7 downto 0);
    signal pc_894 : std_logic_vector(7 downto 0);
    signal type_cast_897_wire_constant : std_logic_vector(7 downto 0);
    signal xxtry1xxzero8 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_zero8_929_wire_constant <= "00000000";
    type_cast_897_wire_constant <= "00000000";
    xxtry1xxzero8 <= "00000000";
    phi_stmt_894: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_897_wire_constant & next_pc_924_898_buffered;
      req <= phi_stmt_894_req_0 & phi_stmt_894_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_894",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_894_ack_0,
          idata => idata,
          odata => pc_894,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_894
    next_pc_924_898_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_pc_924_898_buf_req_0;
      next_pc_924_898_buf_ack_0<= wack(0);
      rreq(0) <= next_pc_924_898_buf_req_1;
      next_pc_924_898_buf_ack_1<= rack(0);
      next_pc_924_898_buf : InterlockBuffer generic map ( -- 
        name => "next_pc_924_898_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_pc_924,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_pc_924_898_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- shared split operator group (0) : CONCAT_u16_u32_919_inst 
    ApConcat_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u8_u16_915_wire & CONCAT_u8_u16_918_wire;
      inst_920 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u16_u32_919_inst_req_0;
      CONCAT_u16_u32_919_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u16_u32_919_inst_req_1;
      CONCAT_u16_u32_919_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_0_gI: SplitGuardInterface generic map(name => "ApConcat_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator CONCAT_u8_u16_915_inst
    process(inst1_902, inst2_905) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(inst1_902, inst2_905, tmp_var);
      CONCAT_u8_u16_915_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_918_inst
    process(inst3_908, inst4_911) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(inst3_908, inst4_911, tmp_var);
      CONCAT_u8_u16_918_wire <= tmp_var; --
    end process;
    -- shared split operator group (3) : CONCAT_u8_u16_931_inst 
    ApConcat_group_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_zero8_929_wire_constant & pc_894;
      CONCAT_u8_u16_931_wire <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u8_u16_931_inst_req_0;
      CONCAT_u8_u16_931_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u8_u16_931_inst_req_1;
      CONCAT_u8_u16_931_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_3_gI: SplitGuardInterface generic map(name => "ApConcat_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared inport operator group (0) : RPIPE_write_mem_904_inst RPIPE_write_mem_910_inst RPIPE_write_mem_907_inst RPIPE_write_mem_901_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 3 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      reqL_unguarded(3) <= RPIPE_write_mem_904_inst_req_0;
      reqL_unguarded(2) <= RPIPE_write_mem_910_inst_req_0;
      reqL_unguarded(1) <= RPIPE_write_mem_907_inst_req_0;
      reqL_unguarded(0) <= RPIPE_write_mem_901_inst_req_0;
      RPIPE_write_mem_904_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_write_mem_910_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_write_mem_907_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_write_mem_901_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= RPIPE_write_mem_904_inst_req_1;
      reqR_unguarded(2) <= RPIPE_write_mem_910_inst_req_1;
      reqR_unguarded(1) <= RPIPE_write_mem_907_inst_req_1;
      reqR_unguarded(0) <= RPIPE_write_mem_901_inst_req_1;
      RPIPE_write_mem_904_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_write_mem_910_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_write_mem_907_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_write_mem_901_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      inst2_905 <= data_out(31 downto 24);
      inst4_911 <= data_out(23 downto 16);
      inst3_908 <= data_out(15 downto 8);
      inst1_902 <= data_out(7 downto 0);
      write_mem_read_0_gI: SplitGuardInterface generic map(name => "write_mem_read_0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      write_mem_read_0: InputPortRevised -- 
        generic map ( name => "write_mem_read_0", data_width => 8,  num_reqs => 4,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => write_mem_pipe_read_req(0),
          oack => write_mem_pipe_read_ack(0),
          odata => write_mem_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_LEDS_928_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LEDS_928_inst_req_0;
      WPIPE_LEDS_928_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LEDS_928_inst_req_1;
      WPIPE_LEDS_928_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= CONCAT_u8_u16_931_wire;
      LEDS_write_0_gI: SplitGuardInterface generic map(name => "LEDS_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LEDS_write_0: OutputPortRevised -- 
        generic map ( name => "LEDS", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LEDS_pipe_write_req(0),
          oack => LEDS_pipe_write_ack(0),
          odata => LEDS_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_reg_output_925_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_reg_output_925_inst_req_0;
      WPIPE_reg_output_925_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_reg_output_925_inst_req_1;
      WPIPE_reg_output_925_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= pc_894;
      reg_output_write_1_gI: SplitGuardInterface generic map(name => "reg_output_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      reg_output_write_1: OutputPortRevised -- 
        generic map ( name => "reg_output", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => reg_output_pipe_write_req(0),
          oack => reg_output_pipe_write_ack(0),
          odata => reg_output_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_890_call 
    init_mem_call_group_0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_890_call_req_0;
      call_stmt_890_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_890_call_req_1;
      call_stmt_890_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      init_mem_call_group_0_gI: SplitGuardInterface generic map(name => "init_mem_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => init_mem_call_reqs(0),
          ackR => init_mem_call_acks(0),
          tagR => init_mem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => init_mem_return_acks(0), -- cross-over
          ackL => init_mem_return_reqs(0), -- cross-over
          tagL => init_mem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_891_call 
    init_reg_call_group_1: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_891_call_req_0;
      call_stmt_891_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_891_call_req_1;
      call_stmt_891_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      init_reg_call_group_1_gI: SplitGuardInterface generic map(name => "init_reg_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => init_reg_call_reqs(0),
          ackR => init_reg_call_acks(0),
          tagR => init_reg_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => init_reg_return_acks(0), -- cross-over
          ackL => init_reg_return_reqs(0), -- cross-over
          tagL => init_reg_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_924_call 
    try_call_group_2: Block -- 
      signal data_in: std_logic_vector(39 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_924_call_req_0;
      call_stmt_924_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_924_call_req_1;
      call_stmt_924_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      try_call_group_2_gI: SplitGuardInterface generic map(name => "try_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= pc_894 & inst_920;
      next_pc_924 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 40,
        owidth => 40,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => try_call_reqs(0),
          ackR => try_call_acks(0),
          dataR => try_call_data(39 downto 0),
          tagR => try_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => try_return_acks(0), -- cross-over
          ackL => try_return_reqs(0), -- cross-over
          dataL => try_return_data(7 downto 0),
          tagL => try_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end try1_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity xnor_i is -- 
  generic (tag_length : integer); 
  port ( -- 
    rs1_data : in  std_logic_vector(31 downto 0);
    rs2_data : in  std_logic_vector(31 downto 0);
    rd : in  std_logic_vector(7 downto 0);
    pc : in  std_logic_vector(7 downto 0);
    next_pc : out  std_logic_vector(7 downto 0);
    accessreg_call_reqs : out  std_logic_vector(0 downto 0);
    accessreg_call_acks : in   std_logic_vector(0 downto 0);
    accessreg_call_data : out  std_logic_vector(40 downto 0);
    accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
    accessreg_return_reqs : out  std_logic_vector(0 downto 0);
    accessreg_return_acks : in   std_logic_vector(0 downto 0);
    accessreg_return_data : in   std_logic_vector(31 downto 0);
    accessreg_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity xnor_i;
architecture xnor_i_arch of xnor_i is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 80)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rs1_data_buffer :  std_logic_vector(31 downto 0);
  signal rs1_data_update_enable: Boolean;
  signal rs2_data_buffer :  std_logic_vector(31 downto 0);
  signal rs2_data_update_enable: Boolean;
  signal rd_buffer :  std_logic_vector(7 downto 0);
  signal rd_update_enable: Boolean;
  signal pc_buffer :  std_logic_vector(7 downto 0);
  signal pc_update_enable: Boolean;
  -- output port buffer signals
  signal next_pc_buffer :  std_logic_vector(7 downto 0);
  signal next_pc_update_enable: Boolean;
  signal xnor_i_CP_1876_start: Boolean;
  signal xnor_i_CP_1876_symbol: Boolean;
  -- volatile/operator module components. 
  component accessreg is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(7 downto 0);
      write_data : in  std_logic_vector(31 downto 0);
      read_data : out  std_logic_vector(31 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal XOR_u32_u32_518_inst_req_0 : boolean;
  signal XOR_u32_u32_518_inst_ack_1 : boolean;
  signal ADD_u8_u8_528_inst_ack_1 : boolean;
  signal call_stmt_524_call_ack_1 : boolean;
  signal XOR_u32_u32_518_inst_req_1 : boolean;
  signal call_stmt_524_call_req_1 : boolean;
  signal call_stmt_524_call_req_0 : boolean;
  signal XOR_u32_u32_518_inst_ack_0 : boolean;
  signal call_stmt_524_call_ack_0 : boolean;
  signal ADD_u8_u8_528_inst_ack_0 : boolean;
  signal ADD_u8_u8_528_inst_req_0 : boolean;
  signal ADD_u8_u8_528_inst_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "xnor_i_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 80) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= rs1_data;
  rs1_data_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= rs2_data;
  rs2_data_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(71 downto 64) <= rd;
  rd_buffer <= in_buffer_data_out(71 downto 64);
  in_buffer_data_in(79 downto 72) <= pc;
  pc_buffer <= in_buffer_data_out(79 downto 72);
  in_buffer_data_in(tag_length + 79 downto 80) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 79 downto 80);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  xnor_i_CP_1876_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "xnor_i_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= next_pc_buffer;
  next_pc <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= xnor_i_CP_1876_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= xnor_i_CP_1876_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= xnor_i_CP_1876_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  xnor_i_CP_1876: Block -- control-path 
    signal xnor_i_CP_1876_elements: BooleanArray(7 downto 0);
    -- 
  begin -- 
    xnor_i_CP_1876_elements(0) <= xnor_i_CP_1876_start;
    xnor_i_CP_1876_symbol <= xnor_i_CP_1876_elements(7);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0:  members (17) 
      -- CP-element group 0: 	 assign_stmt_519_to_assign_stmt_529/call_stmt_524_Update/$entry
      -- CP-element group 0: 	 assign_stmt_519_to_assign_stmt_529/XOR_u32_u32_518_Sample/rr
      -- CP-element group 0: 	 assign_stmt_519_to_assign_stmt_529/ADD_u8_u8_528_sample_start_
      -- CP-element group 0: 	 assign_stmt_519_to_assign_stmt_529/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_519_to_assign_stmt_529/XOR_u32_u32_518_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_519_to_assign_stmt_529/ADD_u8_u8_528_update_start_
      -- CP-element group 0: 	 assign_stmt_519_to_assign_stmt_529/ADD_u8_u8_528_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_519_to_assign_stmt_529/XOR_u32_u32_518_update_start_
      -- CP-element group 0: 	 assign_stmt_519_to_assign_stmt_529/call_stmt_524_update_start_
      -- CP-element group 0: 	 assign_stmt_519_to_assign_stmt_529/XOR_u32_u32_518_sample_start_
      -- CP-element group 0: 	 assign_stmt_519_to_assign_stmt_529/XOR_u32_u32_518_Update/$entry
      -- CP-element group 0: 	 assign_stmt_519_to_assign_stmt_529/XOR_u32_u32_518_Update/cr
      -- CP-element group 0: 	 assign_stmt_519_to_assign_stmt_529/call_stmt_524_Update/ccr
      -- CP-element group 0: 	 assign_stmt_519_to_assign_stmt_529/ADD_u8_u8_528_Update/$entry
      -- CP-element group 0: 	 assign_stmt_519_to_assign_stmt_529/ADD_u8_u8_528_Sample/rr
      -- CP-element group 0: 	 assign_stmt_519_to_assign_stmt_529/ADD_u8_u8_528_Update/cr
      -- 
    cr_1894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => xnor_i_CP_1876_elements(0), ack => XOR_u32_u32_518_inst_req_1); -- 
    ccr_1908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => xnor_i_CP_1876_elements(0), ack => call_stmt_524_call_req_1); -- 
    rr_1917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => xnor_i_CP_1876_elements(0), ack => ADD_u8_u8_528_inst_req_0); -- 
    cr_1922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => xnor_i_CP_1876_elements(0), ack => ADD_u8_u8_528_inst_req_1); -- 
    rr_1889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => xnor_i_CP_1876_elements(0), ack => XOR_u32_u32_518_inst_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_519_to_assign_stmt_529/XOR_u32_u32_518_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_519_to_assign_stmt_529/XOR_u32_u32_518_Sample/ra
      -- CP-element group 1: 	 assign_stmt_519_to_assign_stmt_529/XOR_u32_u32_518_sample_completed_
      -- 
    ra_1890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u32_u32_518_inst_ack_0, ack => xnor_i_CP_1876_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_519_to_assign_stmt_529/call_stmt_524_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_519_to_assign_stmt_529/XOR_u32_u32_518_Update/ca
      -- CP-element group 2: 	 assign_stmt_519_to_assign_stmt_529/XOR_u32_u32_518_Update/$exit
      -- CP-element group 2: 	 assign_stmt_519_to_assign_stmt_529/call_stmt_524_sample_start_
      -- CP-element group 2: 	 assign_stmt_519_to_assign_stmt_529/XOR_u32_u32_518_update_completed_
      -- CP-element group 2: 	 assign_stmt_519_to_assign_stmt_529/call_stmt_524_Sample/crr
      -- 
    ca_1895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u32_u32_518_inst_ack_1, ack => xnor_i_CP_1876_elements(2)); -- 
    crr_1903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => xnor_i_CP_1876_elements(2), ack => call_stmt_524_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_519_to_assign_stmt_529/call_stmt_524_sample_completed_
      -- CP-element group 3: 	 assign_stmt_519_to_assign_stmt_529/call_stmt_524_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_519_to_assign_stmt_529/call_stmt_524_Sample/cra
      -- 
    cra_1904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_524_call_ack_0, ack => xnor_i_CP_1876_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_519_to_assign_stmt_529/call_stmt_524_Update/cca
      -- CP-element group 4: 	 assign_stmt_519_to_assign_stmt_529/call_stmt_524_Update/$exit
      -- CP-element group 4: 	 assign_stmt_519_to_assign_stmt_529/call_stmt_524_update_completed_
      -- 
    cca_1909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_524_call_ack_1, ack => xnor_i_CP_1876_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_519_to_assign_stmt_529/ADD_u8_u8_528_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_519_to_assign_stmt_529/ADD_u8_u8_528_Sample/ra
      -- CP-element group 5: 	 assign_stmt_519_to_assign_stmt_529/ADD_u8_u8_528_sample_completed_
      -- 
    ra_1918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_528_inst_ack_0, ack => xnor_i_CP_1876_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_519_to_assign_stmt_529/ADD_u8_u8_528_Update/ca
      -- CP-element group 6: 	 assign_stmt_519_to_assign_stmt_529/ADD_u8_u8_528_update_completed_
      -- CP-element group 6: 	 assign_stmt_519_to_assign_stmt_529/ADD_u8_u8_528_Update/$exit
      -- 
    ca_1923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_528_inst_ack_1, ack => xnor_i_CP_1876_elements(6)); -- 
    -- CP-element group 7:  join  transition  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 assign_stmt_519_to_assign_stmt_529/$exit
      -- CP-element group 7: 	 $exit
      -- 
    xnor_i_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "xnor_i_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= xnor_i_CP_1876_elements(4) & xnor_i_CP_1876_elements(6);
      gj_xnor_i_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => xnor_i_CP_1876_elements(7), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal dummy_524 : std_logic_vector(31 downto 0);
    signal konst_520_wire_constant : std_logic_vector(0 downto 0);
    signal konst_527_wire_constant : std_logic_vector(7 downto 0);
    signal output_519 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_520_wire_constant <= "0";
    konst_527_wire_constant <= "00000001";
    -- shared split operator group (0) : ADD_u8_u8_528_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pc_buffer;
      next_pc_buffer <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_528_inst_req_0;
      ADD_u8_u8_528_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_528_inst_req_1;
      ADD_u8_u8_528_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : XOR_u32_u32_518_inst 
    ApIntXnor_group_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= rs1_data_buffer & rs2_data_buffer;
      output_519 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= XOR_u32_u32_518_inst_req_0;
      XOR_u32_u32_518_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= XOR_u32_u32_518_inst_req_1;
      XOR_u32_u32_518_inst_ack_1 <= ackR_unguarded(0);
      ApIntXnor_group_1_gI: SplitGuardInterface generic map(name => "ApIntXnor_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntXnor",
          name => "ApIntXnor_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared call operator group (0) : call_stmt_524_call 
    accessreg_call_group_0: Block -- 
      signal data_in: std_logic_vector(40 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_524_call_req_0;
      call_stmt_524_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_524_call_req_1;
      call_stmt_524_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessreg_call_group_0_gI: SplitGuardInterface generic map(name => "accessreg_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_520_wire_constant & rd_buffer & output_519;
      dummy_524 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 41,
        owidth => 41,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessreg_call_reqs(0),
          ackR => accessreg_call_acks(0),
          dataR => accessreg_call_data(40 downto 0),
          tagR => accessreg_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessreg_return_acks(0), -- cross-over
          ackL => accessreg_return_reqs(0), -- cross-over
          dataL => accessreg_return_data(31 downto 0),
          tagL => accessreg_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end xnor_i_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity xor_i is -- 
  generic (tag_length : integer); 
  port ( -- 
    rs1_data : in  std_logic_vector(31 downto 0);
    rs2_data : in  std_logic_vector(31 downto 0);
    rd : in  std_logic_vector(7 downto 0);
    pc : in  std_logic_vector(7 downto 0);
    next_pc : out  std_logic_vector(7 downto 0);
    accessreg_call_reqs : out  std_logic_vector(0 downto 0);
    accessreg_call_acks : in   std_logic_vector(0 downto 0);
    accessreg_call_data : out  std_logic_vector(40 downto 0);
    accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
    accessreg_return_reqs : out  std_logic_vector(0 downto 0);
    accessreg_return_acks : in   std_logic_vector(0 downto 0);
    accessreg_return_data : in   std_logic_vector(31 downto 0);
    accessreg_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity xor_i;
architecture xor_i_arch of xor_i is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 80)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rs1_data_buffer :  std_logic_vector(31 downto 0);
  signal rs1_data_update_enable: Boolean;
  signal rs2_data_buffer :  std_logic_vector(31 downto 0);
  signal rs2_data_update_enable: Boolean;
  signal rd_buffer :  std_logic_vector(7 downto 0);
  signal rd_update_enable: Boolean;
  signal pc_buffer :  std_logic_vector(7 downto 0);
  signal pc_update_enable: Boolean;
  -- output port buffer signals
  signal next_pc_buffer :  std_logic_vector(7 downto 0);
  signal next_pc_update_enable: Boolean;
  signal xor_i_CP_1924_start: Boolean;
  signal xor_i_CP_1924_symbol: Boolean;
  -- volatile/operator module components. 
  component accessreg is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(7 downto 0);
      write_data : in  std_logic_vector(31 downto 0);
      read_data : out  std_logic_vector(31 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal XOR_u32_u32_540_inst_req_0 : boolean;
  signal XOR_u32_u32_540_inst_ack_0 : boolean;
  signal XOR_u32_u32_540_inst_req_1 : boolean;
  signal XOR_u32_u32_540_inst_ack_1 : boolean;
  signal call_stmt_546_call_req_0 : boolean;
  signal call_stmt_546_call_ack_0 : boolean;
  signal call_stmt_546_call_req_1 : boolean;
  signal call_stmt_546_call_ack_1 : boolean;
  signal ADD_u8_u8_550_inst_req_0 : boolean;
  signal ADD_u8_u8_550_inst_ack_0 : boolean;
  signal ADD_u8_u8_550_inst_req_1 : boolean;
  signal ADD_u8_u8_550_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "xor_i_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 80) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= rs1_data;
  rs1_data_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= rs2_data;
  rs2_data_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(71 downto 64) <= rd;
  rd_buffer <= in_buffer_data_out(71 downto 64);
  in_buffer_data_in(79 downto 72) <= pc;
  pc_buffer <= in_buffer_data_out(79 downto 72);
  in_buffer_data_in(tag_length + 79 downto 80) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 79 downto 80);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  xor_i_CP_1924_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "xor_i_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= next_pc_buffer;
  next_pc <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= xor_i_CP_1924_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= xor_i_CP_1924_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= xor_i_CP_1924_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  xor_i_CP_1924: Block -- control-path 
    signal xor_i_CP_1924_elements: BooleanArray(7 downto 0);
    -- 
  begin -- 
    xor_i_CP_1924_elements(0) <= xor_i_CP_1924_start;
    xor_i_CP_1924_symbol <= xor_i_CP_1924_elements(7);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0:  members (17) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_541_to_assign_stmt_551/$entry
      -- CP-element group 0: 	 assign_stmt_541_to_assign_stmt_551/XOR_u32_u32_540_sample_start_
      -- CP-element group 0: 	 assign_stmt_541_to_assign_stmt_551/XOR_u32_u32_540_update_start_
      -- CP-element group 0: 	 assign_stmt_541_to_assign_stmt_551/XOR_u32_u32_540_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_541_to_assign_stmt_551/XOR_u32_u32_540_Sample/rr
      -- CP-element group 0: 	 assign_stmt_541_to_assign_stmt_551/XOR_u32_u32_540_Update/$entry
      -- CP-element group 0: 	 assign_stmt_541_to_assign_stmt_551/XOR_u32_u32_540_Update/cr
      -- CP-element group 0: 	 assign_stmt_541_to_assign_stmt_551/call_stmt_546_update_start_
      -- CP-element group 0: 	 assign_stmt_541_to_assign_stmt_551/call_stmt_546_Update/$entry
      -- CP-element group 0: 	 assign_stmt_541_to_assign_stmt_551/call_stmt_546_Update/ccr
      -- CP-element group 0: 	 assign_stmt_541_to_assign_stmt_551/ADD_u8_u8_550_sample_start_
      -- CP-element group 0: 	 assign_stmt_541_to_assign_stmt_551/ADD_u8_u8_550_update_start_
      -- CP-element group 0: 	 assign_stmt_541_to_assign_stmt_551/ADD_u8_u8_550_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_541_to_assign_stmt_551/ADD_u8_u8_550_Sample/rr
      -- CP-element group 0: 	 assign_stmt_541_to_assign_stmt_551/ADD_u8_u8_550_Update/$entry
      -- CP-element group 0: 	 assign_stmt_541_to_assign_stmt_551/ADD_u8_u8_550_Update/cr
      -- 
    cr_1942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => xor_i_CP_1924_elements(0), ack => XOR_u32_u32_540_inst_req_1); -- 
    rr_1937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => xor_i_CP_1924_elements(0), ack => XOR_u32_u32_540_inst_req_0); -- 
    ccr_1956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => xor_i_CP_1924_elements(0), ack => call_stmt_546_call_req_1); -- 
    rr_1965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => xor_i_CP_1924_elements(0), ack => ADD_u8_u8_550_inst_req_0); -- 
    cr_1970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => xor_i_CP_1924_elements(0), ack => ADD_u8_u8_550_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_541_to_assign_stmt_551/XOR_u32_u32_540_sample_completed_
      -- CP-element group 1: 	 assign_stmt_541_to_assign_stmt_551/XOR_u32_u32_540_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_541_to_assign_stmt_551/XOR_u32_u32_540_Sample/ra
      -- 
    ra_1938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u32_u32_540_inst_ack_0, ack => xor_i_CP_1924_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_541_to_assign_stmt_551/XOR_u32_u32_540_update_completed_
      -- CP-element group 2: 	 assign_stmt_541_to_assign_stmt_551/XOR_u32_u32_540_Update/$exit
      -- CP-element group 2: 	 assign_stmt_541_to_assign_stmt_551/XOR_u32_u32_540_Update/ca
      -- CP-element group 2: 	 assign_stmt_541_to_assign_stmt_551/call_stmt_546_sample_start_
      -- CP-element group 2: 	 assign_stmt_541_to_assign_stmt_551/call_stmt_546_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_541_to_assign_stmt_551/call_stmt_546_Sample/crr
      -- 
    ca_1943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => XOR_u32_u32_540_inst_ack_1, ack => xor_i_CP_1924_elements(2)); -- 
    crr_1951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => xor_i_CP_1924_elements(2), ack => call_stmt_546_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_541_to_assign_stmt_551/call_stmt_546_sample_completed_
      -- CP-element group 3: 	 assign_stmt_541_to_assign_stmt_551/call_stmt_546_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_541_to_assign_stmt_551/call_stmt_546_Sample/cra
      -- 
    cra_1952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_546_call_ack_0, ack => xor_i_CP_1924_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_541_to_assign_stmt_551/call_stmt_546_update_completed_
      -- CP-element group 4: 	 assign_stmt_541_to_assign_stmt_551/call_stmt_546_Update/$exit
      -- CP-element group 4: 	 assign_stmt_541_to_assign_stmt_551/call_stmt_546_Update/cca
      -- 
    cca_1957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_546_call_ack_1, ack => xor_i_CP_1924_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_541_to_assign_stmt_551/ADD_u8_u8_550_sample_completed_
      -- CP-element group 5: 	 assign_stmt_541_to_assign_stmt_551/ADD_u8_u8_550_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_541_to_assign_stmt_551/ADD_u8_u8_550_Sample/ra
      -- 
    ra_1966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_550_inst_ack_0, ack => xor_i_CP_1924_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_541_to_assign_stmt_551/ADD_u8_u8_550_update_completed_
      -- CP-element group 6: 	 assign_stmt_541_to_assign_stmt_551/ADD_u8_u8_550_Update/$exit
      -- CP-element group 6: 	 assign_stmt_541_to_assign_stmt_551/ADD_u8_u8_550_Update/ca
      -- 
    ca_1971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_550_inst_ack_1, ack => xor_i_CP_1924_elements(6)); -- 
    -- CP-element group 7:  join  transition  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 $exit
      -- CP-element group 7: 	 assign_stmt_541_to_assign_stmt_551/$exit
      -- 
    xor_i_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "xor_i_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= xor_i_CP_1924_elements(4) & xor_i_CP_1924_elements(6);
      gj_xor_i_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => xor_i_CP_1924_elements(7), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal dummy_546 : std_logic_vector(31 downto 0);
    signal konst_542_wire_constant : std_logic_vector(0 downto 0);
    signal konst_549_wire_constant : std_logic_vector(7 downto 0);
    signal output_541 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_542_wire_constant <= "0";
    konst_549_wire_constant <= "00000001";
    -- shared split operator group (0) : ADD_u8_u8_550_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pc_buffer;
      next_pc_buffer <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_550_inst_req_0;
      ADD_u8_u8_550_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_550_inst_req_1;
      ADD_u8_u8_550_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : XOR_u32_u32_540_inst 
    ApIntXor_group_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= rs1_data_buffer & rs2_data_buffer;
      output_541 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= XOR_u32_u32_540_inst_req_0;
      XOR_u32_u32_540_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= XOR_u32_u32_540_inst_req_1;
      XOR_u32_u32_540_inst_ack_1 <= ackR_unguarded(0);
      ApIntXor_group_1_gI: SplitGuardInterface generic map(name => "ApIntXor_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          name => "ApIntXor_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared call operator group (0) : call_stmt_546_call 
    accessreg_call_group_0: Block -- 
      signal data_in: std_logic_vector(40 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_546_call_req_0;
      call_stmt_546_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_546_call_req_1;
      call_stmt_546_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessreg_call_group_0_gI: SplitGuardInterface generic map(name => "accessreg_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= konst_542_wire_constant & rd_buffer & output_541;
      dummy_546 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 41,
        owidth => 41,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessreg_call_reqs(0),
          ackR => accessreg_call_acks(0),
          dataR => accessreg_call_data(40 downto 0),
          tagR => accessreg_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessreg_return_acks(0), -- cross-over
          ackL => accessreg_return_reqs(0), -- cross-over
          dataL => accessreg_return_data(31 downto 0),
          tagL => accessreg_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end xor_i_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    LEDS: out std_logic_vector(15 downto 0);
    reg_output_pipe_read_data: out std_logic_vector(7 downto 0);
    reg_output_pipe_read_req : in std_logic_vector(0 downto 0);
    reg_output_pipe_read_ack : out std_logic_vector(0 downto 0);
    write_mem_pipe_write_data: in std_logic_vector(7 downto 0);
    write_mem_pipe_write_req : in std_logic_vector(0 downto 0);
    write_mem_pipe_write_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(7 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(15 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(35 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(2 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(2 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(2 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(59 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(2 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(2 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(23 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(5 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(2 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(2 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(2 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(23 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(59 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(2 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(2 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(5 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(7 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(15 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(35 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(2 downto 0);
  -- declarations related to module accessMem
  component accessMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(7 downto 0);
      write_data : in  std_logic_vector(31 downto 0);
      read_data : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessMem
  signal accessMem_read_write_bar :  std_logic_vector(0 downto 0);
  signal accessMem_addr :  std_logic_vector(7 downto 0);
  signal accessMem_write_data :  std_logic_vector(31 downto 0);
  signal accessMem_read_data :  std_logic_vector(31 downto 0);
  signal accessMem_in_args    : std_logic_vector(40 downto 0);
  signal accessMem_out_args   : std_logic_vector(31 downto 0);
  signal accessMem_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal accessMem_tag_out   : std_logic_vector(2 downto 0);
  signal accessMem_start_req : std_logic;
  signal accessMem_start_ack : std_logic;
  signal accessMem_fin_req   : std_logic;
  signal accessMem_fin_ack : std_logic;
  -- caller side aggregated signals for module accessMem
  signal accessMem_call_reqs: std_logic_vector(1 downto 0);
  signal accessMem_call_acks: std_logic_vector(1 downto 0);
  signal accessMem_return_reqs: std_logic_vector(1 downto 0);
  signal accessMem_return_acks: std_logic_vector(1 downto 0);
  signal accessMem_call_data: std_logic_vector(81 downto 0);
  signal accessMem_call_tag: std_logic_vector(1 downto 0);
  signal accessMem_return_data: std_logic_vector(63 downto 0);
  signal accessMem_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module accessreg
  component accessreg is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar : in  std_logic_vector(0 downto 0);
      addr : in  std_logic_vector(7 downto 0);
      write_data : in  std_logic_vector(31 downto 0);
      read_data : out  std_logic_vector(31 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessreg
  signal accessreg_read_write_bar :  std_logic_vector(0 downto 0);
  signal accessreg_addr :  std_logic_vector(7 downto 0);
  signal accessreg_write_data :  std_logic_vector(31 downto 0);
  signal accessreg_read_data :  std_logic_vector(31 downto 0);
  signal accessreg_in_args    : std_logic_vector(40 downto 0);
  signal accessreg_out_args   : std_logic_vector(31 downto 0);
  signal accessreg_tag_in    : std_logic_vector(5 downto 0) := (others => '0');
  signal accessreg_tag_out   : std_logic_vector(5 downto 0);
  signal accessreg_start_req : std_logic;
  signal accessreg_start_ack : std_logic;
  signal accessreg_fin_req   : std_logic;
  signal accessreg_fin_ack : std_logic;
  -- caller side aggregated signals for module accessreg
  signal accessreg_call_reqs: std_logic_vector(13 downto 0);
  signal accessreg_call_acks: std_logic_vector(13 downto 0);
  signal accessreg_return_reqs: std_logic_vector(13 downto 0);
  signal accessreg_return_acks: std_logic_vector(13 downto 0);
  signal accessreg_call_data: std_logic_vector(573 downto 0);
  signal accessreg_call_tag: std_logic_vector(27 downto 0);
  signal accessreg_return_data: std_logic_vector(447 downto 0);
  signal accessreg_return_tag: std_logic_vector(27 downto 0);
  -- declarations related to module add
  component add is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module add
  signal add_rs1_data :  std_logic_vector(31 downto 0);
  signal add_rs2_data :  std_logic_vector(31 downto 0);
  signal add_rd :  std_logic_vector(7 downto 0);
  signal add_pc :  std_logic_vector(7 downto 0);
  signal add_next_pc :  std_logic_vector(7 downto 0);
  signal add_in_args    : std_logic_vector(79 downto 0);
  signal add_out_args   : std_logic_vector(7 downto 0);
  signal add_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal add_tag_out   : std_logic_vector(1 downto 0);
  signal add_start_req : std_logic;
  signal add_start_ack : std_logic;
  signal add_fin_req   : std_logic;
  signal add_fin_ack : std_logic;
  -- caller side aggregated signals for module add
  signal add_call_reqs: std_logic_vector(0 downto 0);
  signal add_call_acks: std_logic_vector(0 downto 0);
  signal add_return_reqs: std_logic_vector(0 downto 0);
  signal add_return_acks: std_logic_vector(0 downto 0);
  signal add_call_data: std_logic_vector(79 downto 0);
  signal add_call_tag: std_logic_vector(0 downto 0);
  signal add_return_data: std_logic_vector(7 downto 0);
  signal add_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module and_i
  component and_i is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module and_i
  signal and_i_rs1_data :  std_logic_vector(31 downto 0);
  signal and_i_rs2_data :  std_logic_vector(31 downto 0);
  signal and_i_rd :  std_logic_vector(7 downto 0);
  signal and_i_pc :  std_logic_vector(7 downto 0);
  signal and_i_next_pc :  std_logic_vector(7 downto 0);
  signal and_i_in_args    : std_logic_vector(79 downto 0);
  signal and_i_out_args   : std_logic_vector(7 downto 0);
  signal and_i_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal and_i_tag_out   : std_logic_vector(1 downto 0);
  signal and_i_start_req : std_logic;
  signal and_i_start_ack : std_logic;
  signal and_i_fin_req   : std_logic;
  signal and_i_fin_ack : std_logic;
  -- caller side aggregated signals for module and_i
  signal and_i_call_reqs: std_logic_vector(0 downto 0);
  signal and_i_call_acks: std_logic_vector(0 downto 0);
  signal and_i_return_reqs: std_logic_vector(0 downto 0);
  signal and_i_return_acks: std_logic_vector(0 downto 0);
  signal and_i_call_data: std_logic_vector(79 downto 0);
  signal and_i_call_tag: std_logic_vector(0 downto 0);
  signal and_i_return_data: std_logic_vector(7 downto 0);
  signal and_i_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module bn
  component bn is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module bn
  signal bn_rs1_data :  std_logic_vector(31 downto 0);
  signal bn_rs2_data :  std_logic_vector(31 downto 0);
  signal bn_rd :  std_logic_vector(7 downto 0);
  signal bn_pc :  std_logic_vector(7 downto 0);
  signal bn_next_pc :  std_logic_vector(7 downto 0);
  signal bn_in_args    : std_logic_vector(79 downto 0);
  signal bn_out_args   : std_logic_vector(7 downto 0);
  signal bn_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal bn_tag_out   : std_logic_vector(1 downto 0);
  signal bn_start_req : std_logic;
  signal bn_start_ack : std_logic;
  signal bn_fin_req   : std_logic;
  signal bn_fin_ack : std_logic;
  -- caller side aggregated signals for module bn
  signal bn_call_reqs: std_logic_vector(0 downto 0);
  signal bn_call_acks: std_logic_vector(0 downto 0);
  signal bn_return_reqs: std_logic_vector(0 downto 0);
  signal bn_return_acks: std_logic_vector(0 downto 0);
  signal bn_call_data: std_logic_vector(79 downto 0);
  signal bn_call_tag: std_logic_vector(0 downto 0);
  signal bn_return_data: std_logic_vector(7 downto 0);
  signal bn_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module bz
  component bz is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module bz
  signal bz_rs1_data :  std_logic_vector(31 downto 0);
  signal bz_rs2_data :  std_logic_vector(31 downto 0);
  signal bz_rd :  std_logic_vector(7 downto 0);
  signal bz_pc :  std_logic_vector(7 downto 0);
  signal bz_next_pc :  std_logic_vector(7 downto 0);
  signal bz_in_args    : std_logic_vector(79 downto 0);
  signal bz_out_args   : std_logic_vector(7 downto 0);
  signal bz_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal bz_tag_out   : std_logic_vector(1 downto 0);
  signal bz_start_req : std_logic;
  signal bz_start_ack : std_logic;
  signal bz_fin_req   : std_logic;
  signal bz_fin_ack : std_logic;
  -- caller side aggregated signals for module bz
  signal bz_call_reqs: std_logic_vector(0 downto 0);
  signal bz_call_acks: std_logic_vector(0 downto 0);
  signal bz_return_reqs: std_logic_vector(0 downto 0);
  signal bz_return_acks: std_logic_vector(0 downto 0);
  signal bz_call_data: std_logic_vector(79 downto 0);
  signal bz_call_tag: std_logic_vector(0 downto 0);
  signal bz_return_data: std_logic_vector(7 downto 0);
  signal bz_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module call
  component call is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module call
  signal call_rs1_data :  std_logic_vector(31 downto 0);
  signal call_rs2_data :  std_logic_vector(31 downto 0);
  signal call_rd :  std_logic_vector(7 downto 0);
  signal call_pc :  std_logic_vector(7 downto 0);
  signal call_next_pc :  std_logic_vector(7 downto 0);
  signal call_in_args    : std_logic_vector(79 downto 0);
  signal call_out_args   : std_logic_vector(7 downto 0);
  signal call_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal call_tag_out   : std_logic_vector(1 downto 0);
  signal call_start_req : std_logic;
  signal call_start_ack : std_logic;
  signal call_fin_req   : std_logic;
  signal call_fin_ack : std_logic;
  -- caller side aggregated signals for module call
  signal call_call_reqs: std_logic_vector(0 downto 0);
  signal call_call_acks: std_logic_vector(0 downto 0);
  signal call_return_reqs: std_logic_vector(0 downto 0);
  signal call_return_acks: std_logic_vector(0 downto 0);
  signal call_call_data: std_logic_vector(79 downto 0);
  signal call_call_tag: std_logic_vector(0 downto 0);
  signal call_return_data: std_logic_vector(7 downto 0);
  signal call_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module cmp
  component cmp is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module cmp
  signal cmp_rs1_data :  std_logic_vector(31 downto 0);
  signal cmp_rs2_data :  std_logic_vector(31 downto 0);
  signal cmp_rd :  std_logic_vector(7 downto 0);
  signal cmp_pc :  std_logic_vector(7 downto 0);
  signal cmp_next_pc :  std_logic_vector(7 downto 0);
  signal cmp_in_args    : std_logic_vector(79 downto 0);
  signal cmp_out_args   : std_logic_vector(7 downto 0);
  signal cmp_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal cmp_tag_out   : std_logic_vector(1 downto 0);
  signal cmp_start_req : std_logic;
  signal cmp_start_ack : std_logic;
  signal cmp_fin_req   : std_logic;
  signal cmp_fin_ack : std_logic;
  -- caller side aggregated signals for module cmp
  signal cmp_call_reqs: std_logic_vector(0 downto 0);
  signal cmp_call_acks: std_logic_vector(0 downto 0);
  signal cmp_return_reqs: std_logic_vector(0 downto 0);
  signal cmp_return_acks: std_logic_vector(0 downto 0);
  signal cmp_call_data: std_logic_vector(79 downto 0);
  signal cmp_call_tag: std_logic_vector(0 downto 0);
  signal cmp_return_data: std_logic_vector(7 downto 0);
  signal cmp_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module halt
  component halt is -- 
    generic (tag_length : integer); 
    port ( -- 
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module halt
  signal halt_pc :  std_logic_vector(7 downto 0);
  signal halt_next_pc :  std_logic_vector(7 downto 0);
  signal halt_in_args    : std_logic_vector(7 downto 0);
  signal halt_out_args   : std_logic_vector(7 downto 0);
  signal halt_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal halt_tag_out   : std_logic_vector(1 downto 0);
  signal halt_start_req : std_logic;
  signal halt_start_ack : std_logic;
  signal halt_fin_req   : std_logic;
  signal halt_fin_ack : std_logic;
  -- caller side aggregated signals for module halt
  signal halt_call_reqs: std_logic_vector(0 downto 0);
  signal halt_call_acks: std_logic_vector(0 downto 0);
  signal halt_return_reqs: std_logic_vector(0 downto 0);
  signal halt_return_acks: std_logic_vector(0 downto 0);
  signal halt_call_data: std_logic_vector(7 downto 0);
  signal halt_call_tag: std_logic_vector(0 downto 0);
  signal halt_return_data: std_logic_vector(7 downto 0);
  signal halt_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module init_mem
  component init_mem is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module init_mem
  signal init_mem_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal init_mem_tag_out   : std_logic_vector(1 downto 0);
  signal init_mem_start_req : std_logic;
  signal init_mem_start_ack : std_logic;
  signal init_mem_fin_req   : std_logic;
  signal init_mem_fin_ack : std_logic;
  -- caller side aggregated signals for module init_mem
  signal init_mem_call_reqs: std_logic_vector(0 downto 0);
  signal init_mem_call_acks: std_logic_vector(0 downto 0);
  signal init_mem_return_reqs: std_logic_vector(0 downto 0);
  signal init_mem_return_acks: std_logic_vector(0 downto 0);
  signal init_mem_call_tag: std_logic_vector(0 downto 0);
  signal init_mem_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module init_reg
  component init_reg is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module init_reg
  signal init_reg_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal init_reg_tag_out   : std_logic_vector(1 downto 0);
  signal init_reg_start_req : std_logic;
  signal init_reg_start_ack : std_logic;
  signal init_reg_fin_req   : std_logic;
  signal init_reg_fin_ack : std_logic;
  -- caller side aggregated signals for module init_reg
  signal init_reg_call_reqs: std_logic_vector(0 downto 0);
  signal init_reg_call_acks: std_logic_vector(0 downto 0);
  signal init_reg_return_reqs: std_logic_vector(0 downto 0);
  signal init_reg_return_acks: std_logic_vector(0 downto 0);
  signal init_reg_call_tag: std_logic_vector(0 downto 0);
  signal init_reg_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module jmp
  component jmp is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module jmp
  signal jmp_rs1_data :  std_logic_vector(31 downto 0);
  signal jmp_pc :  std_logic_vector(7 downto 0);
  signal jmp_next_pc :  std_logic_vector(7 downto 0);
  signal jmp_in_args    : std_logic_vector(39 downto 0);
  signal jmp_out_args   : std_logic_vector(7 downto 0);
  signal jmp_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal jmp_tag_out   : std_logic_vector(1 downto 0);
  signal jmp_start_req : std_logic;
  signal jmp_start_ack : std_logic;
  signal jmp_fin_req   : std_logic;
  signal jmp_fin_ack : std_logic;
  -- caller side aggregated signals for module jmp
  signal jmp_call_reqs: std_logic_vector(0 downto 0);
  signal jmp_call_acks: std_logic_vector(0 downto 0);
  signal jmp_return_reqs: std_logic_vector(0 downto 0);
  signal jmp_return_acks: std_logic_vector(0 downto 0);
  signal jmp_call_data: std_logic_vector(39 downto 0);
  signal jmp_call_tag: std_logic_vector(0 downto 0);
  signal jmp_return_data: std_logic_vector(7 downto 0);
  signal jmp_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module load
  component load is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessMem_call_acks : in   std_logic_vector(0 downto 0);
      accessMem_call_data : out  std_logic_vector(40 downto 0);
      accessMem_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessMem_return_acks : in   std_logic_vector(0 downto 0);
      accessMem_return_data : in   std_logic_vector(31 downto 0);
      accessMem_return_tag :  in   std_logic_vector(0 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module load
  signal load_rs1_data :  std_logic_vector(31 downto 0);
  signal load_rd :  std_logic_vector(7 downto 0);
  signal load_pc :  std_logic_vector(7 downto 0);
  signal load_next_pc :  std_logic_vector(7 downto 0);
  signal load_in_args    : std_logic_vector(47 downto 0);
  signal load_out_args   : std_logic_vector(7 downto 0);
  signal load_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal load_tag_out   : std_logic_vector(1 downto 0);
  signal load_start_req : std_logic;
  signal load_start_ack : std_logic;
  signal load_fin_req   : std_logic;
  signal load_fin_ack : std_logic;
  -- caller side aggregated signals for module load
  signal load_call_reqs: std_logic_vector(0 downto 0);
  signal load_call_acks: std_logic_vector(0 downto 0);
  signal load_return_reqs: std_logic_vector(0 downto 0);
  signal load_return_acks: std_logic_vector(0 downto 0);
  signal load_call_data: std_logic_vector(47 downto 0);
  signal load_call_tag: std_logic_vector(0 downto 0);
  signal load_return_data: std_logic_vector(7 downto 0);
  signal load_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module or_i
  component or_i is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module or_i
  signal or_i_rs1_data :  std_logic_vector(31 downto 0);
  signal or_i_rs2_data :  std_logic_vector(31 downto 0);
  signal or_i_rd :  std_logic_vector(7 downto 0);
  signal or_i_pc :  std_logic_vector(7 downto 0);
  signal or_i_next_pc :  std_logic_vector(7 downto 0);
  signal or_i_in_args    : std_logic_vector(79 downto 0);
  signal or_i_out_args   : std_logic_vector(7 downto 0);
  signal or_i_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal or_i_tag_out   : std_logic_vector(1 downto 0);
  signal or_i_start_req : std_logic;
  signal or_i_start_ack : std_logic;
  signal or_i_fin_req   : std_logic;
  signal or_i_fin_ack : std_logic;
  -- caller side aggregated signals for module or_i
  signal or_i_call_reqs: std_logic_vector(0 downto 0);
  signal or_i_call_acks: std_logic_vector(0 downto 0);
  signal or_i_return_reqs: std_logic_vector(0 downto 0);
  signal or_i_return_acks: std_logic_vector(0 downto 0);
  signal or_i_call_data: std_logic_vector(79 downto 0);
  signal or_i_call_tag: std_logic_vector(0 downto 0);
  signal or_i_return_data: std_logic_vector(7 downto 0);
  signal or_i_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module sbir
  component sbir is -- 
    generic (tag_length : integer); 
    port ( -- 
      imm : in  std_logic_vector(7 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sbir
  signal sbir_imm :  std_logic_vector(7 downto 0);
  signal sbir_rd :  std_logic_vector(7 downto 0);
  signal sbir_pc :  std_logic_vector(7 downto 0);
  signal sbir_next_pc :  std_logic_vector(7 downto 0);
  signal sbir_in_args    : std_logic_vector(23 downto 0);
  signal sbir_out_args   : std_logic_vector(7 downto 0);
  signal sbir_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sbir_tag_out   : std_logic_vector(1 downto 0);
  signal sbir_start_req : std_logic;
  signal sbir_start_ack : std_logic;
  signal sbir_fin_req   : std_logic;
  signal sbir_fin_ack : std_logic;
  -- caller side aggregated signals for module sbir
  signal sbir_call_reqs: std_logic_vector(0 downto 0);
  signal sbir_call_acks: std_logic_vector(0 downto 0);
  signal sbir_return_reqs: std_logic_vector(0 downto 0);
  signal sbir_return_acks: std_logic_vector(0 downto 0);
  signal sbir_call_data: std_logic_vector(23 downto 0);
  signal sbir_call_tag: std_logic_vector(0 downto 0);
  signal sbir_return_data: std_logic_vector(7 downto 0);
  signal sbir_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module sll_i
  component sll_i is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sll_i
  signal sll_i_rs1_data :  std_logic_vector(31 downto 0);
  signal sll_i_rs2_data :  std_logic_vector(31 downto 0);
  signal sll_i_rd :  std_logic_vector(7 downto 0);
  signal sll_i_pc :  std_logic_vector(7 downto 0);
  signal sll_i_next_pc :  std_logic_vector(7 downto 0);
  signal sll_i_in_args    : std_logic_vector(79 downto 0);
  signal sll_i_out_args   : std_logic_vector(7 downto 0);
  signal sll_i_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sll_i_tag_out   : std_logic_vector(1 downto 0);
  signal sll_i_start_req : std_logic;
  signal sll_i_start_ack : std_logic;
  signal sll_i_fin_req   : std_logic;
  signal sll_i_fin_ack : std_logic;
  -- caller side aggregated signals for module sll_i
  signal sll_i_call_reqs: std_logic_vector(0 downto 0);
  signal sll_i_call_acks: std_logic_vector(0 downto 0);
  signal sll_i_return_reqs: std_logic_vector(0 downto 0);
  signal sll_i_return_acks: std_logic_vector(0 downto 0);
  signal sll_i_call_data: std_logic_vector(79 downto 0);
  signal sll_i_call_tag: std_logic_vector(0 downto 0);
  signal sll_i_return_data: std_logic_vector(7 downto 0);
  signal sll_i_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module sra_i
  component sra_i is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(2 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sra_i
  signal sra_i_rs1_data :  std_logic_vector(31 downto 0);
  signal sra_i_rs2_data :  std_logic_vector(31 downto 0);
  signal sra_i_rd :  std_logic_vector(7 downto 0);
  signal sra_i_pc :  std_logic_vector(7 downto 0);
  signal sra_i_next_pc :  std_logic_vector(7 downto 0);
  signal sra_i_in_args    : std_logic_vector(79 downto 0);
  signal sra_i_out_args   : std_logic_vector(7 downto 0);
  signal sra_i_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sra_i_tag_out   : std_logic_vector(1 downto 0);
  signal sra_i_start_req : std_logic;
  signal sra_i_start_ack : std_logic;
  signal sra_i_fin_req   : std_logic;
  signal sra_i_fin_ack : std_logic;
  -- caller side aggregated signals for module sra_i
  signal sra_i_call_reqs: std_logic_vector(0 downto 0);
  signal sra_i_call_acks: std_logic_vector(0 downto 0);
  signal sra_i_return_reqs: std_logic_vector(0 downto 0);
  signal sra_i_return_acks: std_logic_vector(0 downto 0);
  signal sra_i_call_data: std_logic_vector(79 downto 0);
  signal sra_i_call_tag: std_logic_vector(0 downto 0);
  signal sra_i_return_data: std_logic_vector(7 downto 0);
  signal sra_i_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module srl_i
  component srl_i is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module srl_i
  signal srl_i_rs1_data :  std_logic_vector(31 downto 0);
  signal srl_i_rs2_data :  std_logic_vector(31 downto 0);
  signal srl_i_rd :  std_logic_vector(7 downto 0);
  signal srl_i_pc :  std_logic_vector(7 downto 0);
  signal srl_i_next_pc :  std_logic_vector(7 downto 0);
  signal srl_i_in_args    : std_logic_vector(79 downto 0);
  signal srl_i_out_args   : std_logic_vector(7 downto 0);
  signal srl_i_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal srl_i_tag_out   : std_logic_vector(1 downto 0);
  signal srl_i_start_req : std_logic;
  signal srl_i_start_ack : std_logic;
  signal srl_i_fin_req   : std_logic;
  signal srl_i_fin_ack : std_logic;
  -- caller side aggregated signals for module srl_i
  signal srl_i_call_reqs: std_logic_vector(0 downto 0);
  signal srl_i_call_acks: std_logic_vector(0 downto 0);
  signal srl_i_return_reqs: std_logic_vector(0 downto 0);
  signal srl_i_return_acks: std_logic_vector(0 downto 0);
  signal srl_i_call_data: std_logic_vector(79 downto 0);
  signal srl_i_call_tag: std_logic_vector(0 downto 0);
  signal srl_i_return_data: std_logic_vector(7 downto 0);
  signal srl_i_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module store
  component store is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessMem_call_acks : in   std_logic_vector(0 downto 0);
      accessMem_call_data : out  std_logic_vector(40 downto 0);
      accessMem_call_tag  :  out  std_logic_vector(0 downto 0);
      accessMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessMem_return_acks : in   std_logic_vector(0 downto 0);
      accessMem_return_data : in   std_logic_vector(31 downto 0);
      accessMem_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module store
  signal store_rs1_data :  std_logic_vector(31 downto 0);
  signal store_rs2_data :  std_logic_vector(31 downto 0);
  signal store_pc :  std_logic_vector(7 downto 0);
  signal store_next_pc :  std_logic_vector(7 downto 0);
  signal store_in_args    : std_logic_vector(71 downto 0);
  signal store_out_args   : std_logic_vector(7 downto 0);
  signal store_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal store_tag_out   : std_logic_vector(1 downto 0);
  signal store_start_req : std_logic;
  signal store_start_ack : std_logic;
  signal store_fin_req   : std_logic;
  signal store_fin_ack : std_logic;
  -- caller side aggregated signals for module store
  signal store_call_reqs: std_logic_vector(0 downto 0);
  signal store_call_acks: std_logic_vector(0 downto 0);
  signal store_return_reqs: std_logic_vector(0 downto 0);
  signal store_return_acks: std_logic_vector(0 downto 0);
  signal store_call_data: std_logic_vector(71 downto 0);
  signal store_call_tag: std_logic_vector(0 downto 0);
  signal store_return_data: std_logic_vector(7 downto 0);
  signal store_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module sub
  component sub is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sub
  signal sub_rs1_data :  std_logic_vector(31 downto 0);
  signal sub_rs2_data :  std_logic_vector(31 downto 0);
  signal sub_rd :  std_logic_vector(7 downto 0);
  signal sub_pc :  std_logic_vector(7 downto 0);
  signal sub_next_pc :  std_logic_vector(7 downto 0);
  signal sub_in_args    : std_logic_vector(79 downto 0);
  signal sub_out_args   : std_logic_vector(7 downto 0);
  signal sub_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sub_tag_out   : std_logic_vector(1 downto 0);
  signal sub_start_req : std_logic;
  signal sub_start_ack : std_logic;
  signal sub_fin_req   : std_logic;
  signal sub_fin_ack : std_logic;
  -- caller side aggregated signals for module sub
  signal sub_call_reqs: std_logic_vector(0 downto 0);
  signal sub_call_acks: std_logic_vector(0 downto 0);
  signal sub_return_reqs: std_logic_vector(0 downto 0);
  signal sub_return_acks: std_logic_vector(0 downto 0);
  signal sub_call_data: std_logic_vector(79 downto 0);
  signal sub_call_tag: std_logic_vector(0 downto 0);
  signal sub_return_data: std_logic_vector(7 downto 0);
  signal sub_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module try
  component try is -- 
    generic (tag_length : integer); 
    port ( -- 
      pc : in  std_logic_vector(7 downto 0);
      inst : in  std_logic_vector(31 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      cmp_call_reqs : out  std_logic_vector(0 downto 0);
      cmp_call_acks : in   std_logic_vector(0 downto 0);
      cmp_call_data : out  std_logic_vector(79 downto 0);
      cmp_call_tag  :  out  std_logic_vector(0 downto 0);
      cmp_return_reqs : out  std_logic_vector(0 downto 0);
      cmp_return_acks : in   std_logic_vector(0 downto 0);
      cmp_return_data : in   std_logic_vector(7 downto 0);
      cmp_return_tag :  in   std_logic_vector(0 downto 0);
      sub_call_reqs : out  std_logic_vector(0 downto 0);
      sub_call_acks : in   std_logic_vector(0 downto 0);
      sub_call_data : out  std_logic_vector(79 downto 0);
      sub_call_tag  :  out  std_logic_vector(0 downto 0);
      sub_return_reqs : out  std_logic_vector(0 downto 0);
      sub_return_acks : in   std_logic_vector(0 downto 0);
      sub_return_data : in   std_logic_vector(7 downto 0);
      sub_return_tag :  in   std_logic_vector(0 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      bn_call_reqs : out  std_logic_vector(0 downto 0);
      bn_call_acks : in   std_logic_vector(0 downto 0);
      bn_call_data : out  std_logic_vector(79 downto 0);
      bn_call_tag  :  out  std_logic_vector(0 downto 0);
      bn_return_reqs : out  std_logic_vector(0 downto 0);
      bn_return_acks : in   std_logic_vector(0 downto 0);
      bn_return_data : in   std_logic_vector(7 downto 0);
      bn_return_tag :  in   std_logic_vector(0 downto 0);
      halt_call_reqs : out  std_logic_vector(0 downto 0);
      halt_call_acks : in   std_logic_vector(0 downto 0);
      halt_call_data : out  std_logic_vector(7 downto 0);
      halt_call_tag  :  out  std_logic_vector(0 downto 0);
      halt_return_reqs : out  std_logic_vector(0 downto 0);
      halt_return_acks : in   std_logic_vector(0 downto 0);
      halt_return_data : in   std_logic_vector(7 downto 0);
      halt_return_tag :  in   std_logic_vector(0 downto 0);
      add_call_reqs : out  std_logic_vector(0 downto 0);
      add_call_acks : in   std_logic_vector(0 downto 0);
      add_call_data : out  std_logic_vector(79 downto 0);
      add_call_tag  :  out  std_logic_vector(0 downto 0);
      add_return_reqs : out  std_logic_vector(0 downto 0);
      add_return_acks : in   std_logic_vector(0 downto 0);
      add_return_data : in   std_logic_vector(7 downto 0);
      add_return_tag :  in   std_logic_vector(0 downto 0);
      sll_i_call_reqs : out  std_logic_vector(0 downto 0);
      sll_i_call_acks : in   std_logic_vector(0 downto 0);
      sll_i_call_data : out  std_logic_vector(79 downto 0);
      sll_i_call_tag  :  out  std_logic_vector(0 downto 0);
      sll_i_return_reqs : out  std_logic_vector(0 downto 0);
      sll_i_return_acks : in   std_logic_vector(0 downto 0);
      sll_i_return_data : in   std_logic_vector(7 downto 0);
      sll_i_return_tag :  in   std_logic_vector(0 downto 0);
      and_i_call_reqs : out  std_logic_vector(0 downto 0);
      and_i_call_acks : in   std_logic_vector(0 downto 0);
      and_i_call_data : out  std_logic_vector(79 downto 0);
      and_i_call_tag  :  out  std_logic_vector(0 downto 0);
      and_i_return_reqs : out  std_logic_vector(0 downto 0);
      and_i_return_acks : in   std_logic_vector(0 downto 0);
      and_i_return_data : in   std_logic_vector(7 downto 0);
      and_i_return_tag :  in   std_logic_vector(0 downto 0);
      call_call_reqs : out  std_logic_vector(0 downto 0);
      call_call_acks : in   std_logic_vector(0 downto 0);
      call_call_data : out  std_logic_vector(79 downto 0);
      call_call_tag  :  out  std_logic_vector(0 downto 0);
      call_return_reqs : out  std_logic_vector(0 downto 0);
      call_return_acks : in   std_logic_vector(0 downto 0);
      call_return_data : in   std_logic_vector(7 downto 0);
      call_return_tag :  in   std_logic_vector(0 downto 0);
      bz_call_reqs : out  std_logic_vector(0 downto 0);
      bz_call_acks : in   std_logic_vector(0 downto 0);
      bz_call_data : out  std_logic_vector(79 downto 0);
      bz_call_tag  :  out  std_logic_vector(0 downto 0);
      bz_return_reqs : out  std_logic_vector(0 downto 0);
      bz_return_acks : in   std_logic_vector(0 downto 0);
      bz_return_data : in   std_logic_vector(7 downto 0);
      bz_return_tag :  in   std_logic_vector(0 downto 0);
      xnor_i_call_reqs : out  std_logic_vector(0 downto 0);
      xnor_i_call_acks : in   std_logic_vector(0 downto 0);
      xnor_i_call_data : out  std_logic_vector(79 downto 0);
      xnor_i_call_tag  :  out  std_logic_vector(0 downto 0);
      xnor_i_return_reqs : out  std_logic_vector(0 downto 0);
      xnor_i_return_acks : in   std_logic_vector(0 downto 0);
      xnor_i_return_data : in   std_logic_vector(7 downto 0);
      xnor_i_return_tag :  in   std_logic_vector(0 downto 0);
      sra_i_call_reqs : out  std_logic_vector(0 downto 0);
      sra_i_call_acks : in   std_logic_vector(0 downto 0);
      sra_i_call_data : out  std_logic_vector(79 downto 0);
      sra_i_call_tag  :  out  std_logic_vector(0 downto 0);
      sra_i_return_reqs : out  std_logic_vector(0 downto 0);
      sra_i_return_acks : in   std_logic_vector(0 downto 0);
      sra_i_return_data : in   std_logic_vector(7 downto 0);
      sra_i_return_tag :  in   std_logic_vector(0 downto 0);
      sbir_call_reqs : out  std_logic_vector(0 downto 0);
      sbir_call_acks : in   std_logic_vector(0 downto 0);
      sbir_call_data : out  std_logic_vector(23 downto 0);
      sbir_call_tag  :  out  std_logic_vector(0 downto 0);
      sbir_return_reqs : out  std_logic_vector(0 downto 0);
      sbir_return_acks : in   std_logic_vector(0 downto 0);
      sbir_return_data : in   std_logic_vector(7 downto 0);
      sbir_return_tag :  in   std_logic_vector(0 downto 0);
      or_i_call_reqs : out  std_logic_vector(0 downto 0);
      or_i_call_acks : in   std_logic_vector(0 downto 0);
      or_i_call_data : out  std_logic_vector(79 downto 0);
      or_i_call_tag  :  out  std_logic_vector(0 downto 0);
      or_i_return_reqs : out  std_logic_vector(0 downto 0);
      or_i_return_acks : in   std_logic_vector(0 downto 0);
      or_i_return_data : in   std_logic_vector(7 downto 0);
      or_i_return_tag :  in   std_logic_vector(0 downto 0);
      load_call_reqs : out  std_logic_vector(0 downto 0);
      load_call_acks : in   std_logic_vector(0 downto 0);
      load_call_data : out  std_logic_vector(47 downto 0);
      load_call_tag  :  out  std_logic_vector(0 downto 0);
      load_return_reqs : out  std_logic_vector(0 downto 0);
      load_return_acks : in   std_logic_vector(0 downto 0);
      load_return_data : in   std_logic_vector(7 downto 0);
      load_return_tag :  in   std_logic_vector(0 downto 0);
      jmp_call_reqs : out  std_logic_vector(0 downto 0);
      jmp_call_acks : in   std_logic_vector(0 downto 0);
      jmp_call_data : out  std_logic_vector(39 downto 0);
      jmp_call_tag  :  out  std_logic_vector(0 downto 0);
      jmp_return_reqs : out  std_logic_vector(0 downto 0);
      jmp_return_acks : in   std_logic_vector(0 downto 0);
      jmp_return_data : in   std_logic_vector(7 downto 0);
      jmp_return_tag :  in   std_logic_vector(0 downto 0);
      store_call_reqs : out  std_logic_vector(0 downto 0);
      store_call_acks : in   std_logic_vector(0 downto 0);
      store_call_data : out  std_logic_vector(71 downto 0);
      store_call_tag  :  out  std_logic_vector(0 downto 0);
      store_return_reqs : out  std_logic_vector(0 downto 0);
      store_return_acks : in   std_logic_vector(0 downto 0);
      store_return_data : in   std_logic_vector(7 downto 0);
      store_return_tag :  in   std_logic_vector(0 downto 0);
      srl_i_call_reqs : out  std_logic_vector(0 downto 0);
      srl_i_call_acks : in   std_logic_vector(0 downto 0);
      srl_i_call_data : out  std_logic_vector(79 downto 0);
      srl_i_call_tag  :  out  std_logic_vector(0 downto 0);
      srl_i_return_reqs : out  std_logic_vector(0 downto 0);
      srl_i_return_acks : in   std_logic_vector(0 downto 0);
      srl_i_return_data : in   std_logic_vector(7 downto 0);
      srl_i_return_tag :  in   std_logic_vector(0 downto 0);
      xor_i_call_reqs : out  std_logic_vector(0 downto 0);
      xor_i_call_acks : in   std_logic_vector(0 downto 0);
      xor_i_call_data : out  std_logic_vector(79 downto 0);
      xor_i_call_tag  :  out  std_logic_vector(0 downto 0);
      xor_i_return_reqs : out  std_logic_vector(0 downto 0);
      xor_i_return_acks : in   std_logic_vector(0 downto 0);
      xor_i_return_data : in   std_logic_vector(7 downto 0);
      xor_i_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module try
  signal try_pc :  std_logic_vector(7 downto 0);
  signal try_inst :  std_logic_vector(31 downto 0);
  signal try_next_pc :  std_logic_vector(7 downto 0);
  signal try_in_args    : std_logic_vector(39 downto 0);
  signal try_out_args   : std_logic_vector(7 downto 0);
  signal try_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal try_tag_out   : std_logic_vector(1 downto 0);
  signal try_start_req : std_logic;
  signal try_start_ack : std_logic;
  signal try_fin_req   : std_logic;
  signal try_fin_ack : std_logic;
  -- caller side aggregated signals for module try
  signal try_call_reqs: std_logic_vector(0 downto 0);
  signal try_call_acks: std_logic_vector(0 downto 0);
  signal try_return_reqs: std_logic_vector(0 downto 0);
  signal try_return_acks: std_logic_vector(0 downto 0);
  signal try_call_data: std_logic_vector(39 downto 0);
  signal try_call_tag: std_logic_vector(0 downto 0);
  signal try_return_data: std_logic_vector(7 downto 0);
  signal try_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module try1
  component try1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      write_mem_pipe_read_req : out  std_logic_vector(0 downto 0);
      write_mem_pipe_read_ack : in   std_logic_vector(0 downto 0);
      write_mem_pipe_read_data : in   std_logic_vector(7 downto 0);
      LEDS_pipe_write_req : out  std_logic_vector(0 downto 0);
      LEDS_pipe_write_ack : in   std_logic_vector(0 downto 0);
      LEDS_pipe_write_data : out  std_logic_vector(15 downto 0);
      reg_output_pipe_write_req : out  std_logic_vector(0 downto 0);
      reg_output_pipe_write_ack : in   std_logic_vector(0 downto 0);
      reg_output_pipe_write_data : out  std_logic_vector(7 downto 0);
      init_mem_call_reqs : out  std_logic_vector(0 downto 0);
      init_mem_call_acks : in   std_logic_vector(0 downto 0);
      init_mem_call_tag  :  out  std_logic_vector(0 downto 0);
      init_mem_return_reqs : out  std_logic_vector(0 downto 0);
      init_mem_return_acks : in   std_logic_vector(0 downto 0);
      init_mem_return_tag :  in   std_logic_vector(0 downto 0);
      init_reg_call_reqs : out  std_logic_vector(0 downto 0);
      init_reg_call_acks : in   std_logic_vector(0 downto 0);
      init_reg_call_tag  :  out  std_logic_vector(0 downto 0);
      init_reg_return_reqs : out  std_logic_vector(0 downto 0);
      init_reg_return_acks : in   std_logic_vector(0 downto 0);
      init_reg_return_tag :  in   std_logic_vector(0 downto 0);
      try_call_reqs : out  std_logic_vector(0 downto 0);
      try_call_acks : in   std_logic_vector(0 downto 0);
      try_call_data : out  std_logic_vector(39 downto 0);
      try_call_tag  :  out  std_logic_vector(0 downto 0);
      try_return_reqs : out  std_logic_vector(0 downto 0);
      try_return_acks : in   std_logic_vector(0 downto 0);
      try_return_data : in   std_logic_vector(7 downto 0);
      try_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module try1
  signal try1_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal try1_tag_out   : std_logic_vector(1 downto 0);
  signal try1_start_req : std_logic;
  signal try1_start_ack : std_logic;
  signal try1_fin_req   : std_logic;
  signal try1_fin_ack : std_logic;
  -- declarations related to module xnor_i
  component xnor_i is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module xnor_i
  signal xnor_i_rs1_data :  std_logic_vector(31 downto 0);
  signal xnor_i_rs2_data :  std_logic_vector(31 downto 0);
  signal xnor_i_rd :  std_logic_vector(7 downto 0);
  signal xnor_i_pc :  std_logic_vector(7 downto 0);
  signal xnor_i_next_pc :  std_logic_vector(7 downto 0);
  signal xnor_i_in_args    : std_logic_vector(79 downto 0);
  signal xnor_i_out_args   : std_logic_vector(7 downto 0);
  signal xnor_i_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal xnor_i_tag_out   : std_logic_vector(1 downto 0);
  signal xnor_i_start_req : std_logic;
  signal xnor_i_start_ack : std_logic;
  signal xnor_i_fin_req   : std_logic;
  signal xnor_i_fin_ack : std_logic;
  -- caller side aggregated signals for module xnor_i
  signal xnor_i_call_reqs: std_logic_vector(0 downto 0);
  signal xnor_i_call_acks: std_logic_vector(0 downto 0);
  signal xnor_i_return_reqs: std_logic_vector(0 downto 0);
  signal xnor_i_return_acks: std_logic_vector(0 downto 0);
  signal xnor_i_call_data: std_logic_vector(79 downto 0);
  signal xnor_i_call_tag: std_logic_vector(0 downto 0);
  signal xnor_i_return_data: std_logic_vector(7 downto 0);
  signal xnor_i_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module xor_i
  component xor_i is -- 
    generic (tag_length : integer); 
    port ( -- 
      rs1_data : in  std_logic_vector(31 downto 0);
      rs2_data : in  std_logic_vector(31 downto 0);
      rd : in  std_logic_vector(7 downto 0);
      pc : in  std_logic_vector(7 downto 0);
      next_pc : out  std_logic_vector(7 downto 0);
      accessreg_call_reqs : out  std_logic_vector(0 downto 0);
      accessreg_call_acks : in   std_logic_vector(0 downto 0);
      accessreg_call_data : out  std_logic_vector(40 downto 0);
      accessreg_call_tag  :  out  std_logic_vector(1 downto 0);
      accessreg_return_reqs : out  std_logic_vector(0 downto 0);
      accessreg_return_acks : in   std_logic_vector(0 downto 0);
      accessreg_return_data : in   std_logic_vector(31 downto 0);
      accessreg_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module xor_i
  signal xor_i_rs1_data :  std_logic_vector(31 downto 0);
  signal xor_i_rs2_data :  std_logic_vector(31 downto 0);
  signal xor_i_rd :  std_logic_vector(7 downto 0);
  signal xor_i_pc :  std_logic_vector(7 downto 0);
  signal xor_i_next_pc :  std_logic_vector(7 downto 0);
  signal xor_i_in_args    : std_logic_vector(79 downto 0);
  signal xor_i_out_args   : std_logic_vector(7 downto 0);
  signal xor_i_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal xor_i_tag_out   : std_logic_vector(1 downto 0);
  signal xor_i_start_req : std_logic;
  signal xor_i_start_ack : std_logic;
  signal xor_i_fin_req   : std_logic;
  signal xor_i_fin_ack : std_logic;
  -- caller side aggregated signals for module xor_i
  signal xor_i_call_reqs: std_logic_vector(0 downto 0);
  signal xor_i_call_acks: std_logic_vector(0 downto 0);
  signal xor_i_return_reqs: std_logic_vector(0 downto 0);
  signal xor_i_return_acks: std_logic_vector(0 downto 0);
  signal xor_i_call_data: std_logic_vector(79 downto 0);
  signal xor_i_call_tag: std_logic_vector(0 downto 0);
  signal xor_i_return_data: std_logic_vector(7 downto 0);
  signal xor_i_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe LEDS
  signal LEDS_pipe_write_data: std_logic_vector(15 downto 0);
  signal LEDS_pipe_write_req: std_logic_vector(0 downto 0);
  signal LEDS_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe reg_output
  signal reg_output_pipe_write_data: std_logic_vector(7 downto 0);
  signal reg_output_pipe_write_req: std_logic_vector(0 downto 0);
  signal reg_output_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe write_mem
  signal write_mem_pipe_read_data: std_logic_vector(7 downto 0);
  signal write_mem_pipe_read_req: std_logic_vector(0 downto 0);
  signal write_mem_pipe_read_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module accessMem
  accessMem_read_write_bar <= accessMem_in_args(40 downto 40);
  accessMem_addr <= accessMem_in_args(39 downto 32);
  accessMem_write_data <= accessMem_in_args(31 downto 0);
  accessMem_out_args <= accessMem_read_data ;
  -- call arbiter for module accessMem
  accessMem_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 41,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => accessMem_call_reqs,
      call_acks => accessMem_call_acks,
      return_reqs => accessMem_return_reqs,
      return_acks => accessMem_return_acks,
      call_data  => accessMem_call_data,
      call_tag  => accessMem_call_tag,
      return_tag  => accessMem_return_tag,
      call_mtag => accessMem_tag_in,
      return_mtag => accessMem_tag_out,
      return_data =>accessMem_return_data,
      call_mreq => accessMem_start_req,
      call_mack => accessMem_start_ack,
      return_mreq => accessMem_fin_req,
      return_mack => accessMem_fin_ack,
      call_mdata => accessMem_in_args,
      return_mdata => accessMem_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessMem_instance:accessMem-- 
    generic map(tag_length => 3)
    port map(-- 
      read_write_bar => accessMem_read_write_bar,
      addr => accessMem_addr,
      write_data => accessMem_write_data,
      read_data => accessMem_read_data,
      start_req => accessMem_start_req,
      start_ack => accessMem_start_ack,
      fin_req => accessMem_fin_req,
      fin_ack => accessMem_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(7 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(17 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(31 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(1 downto 1),
      memory_space_0_sr_ack => memory_space_0_sr_ack(1 downto 1),
      memory_space_0_sr_addr => memory_space_0_sr_addr(15 downto 8),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 32),
      memory_space_0_sr_tag => memory_space_0_sr_tag(35 downto 18),
      memory_space_0_sc_req => memory_space_0_sc_req(1 downto 1),
      memory_space_0_sc_ack => memory_space_0_sc_ack(1 downto 1),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 1),
      tag_in => accessMem_tag_in,
      tag_out => accessMem_tag_out-- 
    ); -- 
  -- module accessreg
  accessreg_read_write_bar <= accessreg_in_args(40 downto 40);
  accessreg_addr <= accessreg_in_args(39 downto 32);
  accessreg_write_data <= accessreg_in_args(31 downto 0);
  accessreg_out_args <= accessreg_read_data ;
  -- call arbiter for module accessreg
  accessreg_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 14,
      call_data_width => 41,
      return_data_width => 32,
      callee_tag_length => 4,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => accessreg_call_reqs,
      call_acks => accessreg_call_acks,
      return_reqs => accessreg_return_reqs,
      return_acks => accessreg_return_acks,
      call_data  => accessreg_call_data,
      call_tag  => accessreg_call_tag,
      return_tag  => accessreg_return_tag,
      call_mtag => accessreg_tag_in,
      return_mtag => accessreg_tag_out,
      return_data =>accessreg_return_data,
      call_mreq => accessreg_start_req,
      call_mack => accessreg_start_ack,
      return_mreq => accessreg_fin_req,
      return_mack => accessreg_fin_ack,
      call_mdata => accessreg_in_args,
      return_mdata => accessreg_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessreg_instance:accessreg-- 
    generic map(tag_length => 6)
    port map(-- 
      read_write_bar => accessreg_read_write_bar,
      addr => accessreg_addr,
      write_data => accessreg_write_data,
      read_data => accessreg_read_data,
      start_req => accessreg_start_req,
      start_ack => accessreg_start_ack,
      fin_req => accessreg_fin_req,
      fin_ack => accessreg_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(7 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(17 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(31 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(1 downto 1),
      memory_space_2_sr_ack => memory_space_2_sr_ack(1 downto 1),
      memory_space_2_sr_addr => memory_space_2_sr_addr(15 downto 8),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 32),
      memory_space_2_sr_tag => memory_space_2_sr_tag(35 downto 18),
      memory_space_2_sc_req => memory_space_2_sc_req(1 downto 1),
      memory_space_2_sc_ack => memory_space_2_sc_ack(1 downto 1),
      memory_space_2_sc_tag => memory_space_2_sc_tag(1 downto 1),
      tag_in => accessreg_tag_in,
      tag_out => accessreg_tag_out-- 
    ); -- 
  -- module add
  add_rs1_data <= add_in_args(79 downto 48);
  add_rs2_data <= add_in_args(47 downto 16);
  add_rd <= add_in_args(15 downto 8);
  add_pc <= add_in_args(7 downto 0);
  add_out_args <= add_next_pc ;
  -- call arbiter for module add
  add_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 80,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => add_call_reqs,
      call_acks => add_call_acks,
      return_reqs => add_return_reqs,
      return_acks => add_return_acks,
      call_data  => add_call_data,
      call_tag  => add_call_tag,
      return_tag  => add_return_tag,
      call_mtag => add_tag_in,
      return_mtag => add_tag_out,
      return_data =>add_return_data,
      call_mreq => add_start_req,
      call_mack => add_start_ack,
      return_mreq => add_fin_req,
      return_mack => add_fin_ack,
      call_mdata => add_in_args,
      return_mdata => add_out_args,
      clk => clk, 
      reset => reset --
    ); --
  add_instance:add-- 
    generic map(tag_length => 2)
    port map(-- 
      rs1_data => add_rs1_data,
      rs2_data => add_rs2_data,
      rd => add_rd,
      pc => add_pc,
      next_pc => add_next_pc,
      start_req => add_start_req,
      start_ack => add_start_ack,
      fin_req => add_fin_req,
      fin_ack => add_fin_ack,
      clk => clk,
      reset => reset,
      accessreg_call_reqs => accessreg_call_reqs(11 downto 11),
      accessreg_call_acks => accessreg_call_acks(11 downto 11),
      accessreg_call_data => accessreg_call_data(491 downto 451),
      accessreg_call_tag => accessreg_call_tag(23 downto 22),
      accessreg_return_reqs => accessreg_return_reqs(11 downto 11),
      accessreg_return_acks => accessreg_return_acks(11 downto 11),
      accessreg_return_data => accessreg_return_data(383 downto 352),
      accessreg_return_tag => accessreg_return_tag(23 downto 22),
      tag_in => add_tag_in,
      tag_out => add_tag_out-- 
    ); -- 
  -- module and_i
  and_i_rs1_data <= and_i_in_args(79 downto 48);
  and_i_rs2_data <= and_i_in_args(47 downto 16);
  and_i_rd <= and_i_in_args(15 downto 8);
  and_i_pc <= and_i_in_args(7 downto 0);
  and_i_out_args <= and_i_next_pc ;
  -- call arbiter for module and_i
  and_i_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 80,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => and_i_call_reqs,
      call_acks => and_i_call_acks,
      return_reqs => and_i_return_reqs,
      return_acks => and_i_return_acks,
      call_data  => and_i_call_data,
      call_tag  => and_i_call_tag,
      return_tag  => and_i_return_tag,
      call_mtag => and_i_tag_in,
      return_mtag => and_i_tag_out,
      return_data =>and_i_return_data,
      call_mreq => and_i_start_req,
      call_mack => and_i_start_ack,
      return_mreq => and_i_fin_req,
      return_mack => and_i_fin_ack,
      call_mdata => and_i_in_args,
      return_mdata => and_i_out_args,
      clk => clk, 
      reset => reset --
    ); --
  and_i_instance:and_i-- 
    generic map(tag_length => 2)
    port map(-- 
      rs1_data => and_i_rs1_data,
      rs2_data => and_i_rs2_data,
      rd => and_i_rd,
      pc => and_i_pc,
      next_pc => and_i_next_pc,
      start_req => and_i_start_req,
      start_ack => and_i_start_ack,
      fin_req => and_i_fin_req,
      fin_ack => and_i_fin_ack,
      clk => clk,
      reset => reset,
      accessreg_call_reqs => accessreg_call_reqs(9 downto 9),
      accessreg_call_acks => accessreg_call_acks(9 downto 9),
      accessreg_call_data => accessreg_call_data(409 downto 369),
      accessreg_call_tag => accessreg_call_tag(19 downto 18),
      accessreg_return_reqs => accessreg_return_reqs(9 downto 9),
      accessreg_return_acks => accessreg_return_acks(9 downto 9),
      accessreg_return_data => accessreg_return_data(319 downto 288),
      accessreg_return_tag => accessreg_return_tag(19 downto 18),
      tag_in => and_i_tag_in,
      tag_out => and_i_tag_out-- 
    ); -- 
  -- module bn
  bn_rs1_data <= bn_in_args(79 downto 48);
  bn_rs2_data <= bn_in_args(47 downto 16);
  bn_rd <= bn_in_args(15 downto 8);
  bn_pc <= bn_in_args(7 downto 0);
  bn_out_args <= bn_next_pc ;
  -- call arbiter for module bn
  bn_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 80,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => bn_call_reqs,
      call_acks => bn_call_acks,
      return_reqs => bn_return_reqs,
      return_acks => bn_return_acks,
      call_data  => bn_call_data,
      call_tag  => bn_call_tag,
      return_tag  => bn_return_tag,
      call_mtag => bn_tag_in,
      return_mtag => bn_tag_out,
      return_data =>bn_return_data,
      call_mreq => bn_start_req,
      call_mack => bn_start_ack,
      return_mreq => bn_fin_req,
      return_mack => bn_fin_ack,
      call_mdata => bn_in_args,
      return_mdata => bn_out_args,
      clk => clk, 
      reset => reset --
    ); --
  bn_instance:bn-- 
    generic map(tag_length => 2)
    port map(-- 
      rs1_data => bn_rs1_data,
      rs2_data => bn_rs2_data,
      rd => bn_rd,
      pc => bn_pc,
      next_pc => bn_next_pc,
      start_req => bn_start_req,
      start_ack => bn_start_ack,
      fin_req => bn_fin_req,
      fin_ack => bn_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(2 downto 2),
      memory_space_1_lr_tag => memory_space_1_lr_tag(59 downto 40),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(23 downto 16),
      memory_space_1_lc_tag => memory_space_1_lc_tag(5 downto 4),
      memory_space_1_sr_req => memory_space_1_sr_req(2 downto 2),
      memory_space_1_sr_ack => memory_space_1_sr_ack(2 downto 2),
      memory_space_1_sr_addr => memory_space_1_sr_addr(2 downto 2),
      memory_space_1_sr_data => memory_space_1_sr_data(23 downto 16),
      memory_space_1_sr_tag => memory_space_1_sr_tag(59 downto 40),
      memory_space_1_sc_req => memory_space_1_sc_req(2 downto 2),
      memory_space_1_sc_ack => memory_space_1_sc_ack(2 downto 2),
      memory_space_1_sc_tag => memory_space_1_sc_tag(5 downto 4),
      tag_in => bn_tag_in,
      tag_out => bn_tag_out-- 
    ); -- 
  -- module bz
  bz_rs1_data <= bz_in_args(79 downto 48);
  bz_rs2_data <= bz_in_args(47 downto 16);
  bz_rd <= bz_in_args(15 downto 8);
  bz_pc <= bz_in_args(7 downto 0);
  bz_out_args <= bz_next_pc ;
  -- call arbiter for module bz
  bz_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 80,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => bz_call_reqs,
      call_acks => bz_call_acks,
      return_reqs => bz_return_reqs,
      return_acks => bz_return_acks,
      call_data  => bz_call_data,
      call_tag  => bz_call_tag,
      return_tag  => bz_return_tag,
      call_mtag => bz_tag_in,
      return_mtag => bz_tag_out,
      return_data =>bz_return_data,
      call_mreq => bz_start_req,
      call_mack => bz_start_ack,
      return_mreq => bz_fin_req,
      return_mack => bz_fin_ack,
      call_mdata => bz_in_args,
      return_mdata => bz_out_args,
      clk => clk, 
      reset => reset --
    ); --
  bz_instance:bz-- 
    generic map(tag_length => 2)
    port map(-- 
      rs1_data => bz_rs1_data,
      rs2_data => bz_rs2_data,
      rd => bz_rd,
      pc => bz_pc,
      next_pc => bz_next_pc,
      start_req => bz_start_req,
      start_ack => bz_start_ack,
      fin_req => bz_fin_req,
      fin_ack => bz_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(1 downto 1),
      memory_space_1_lr_tag => memory_space_1_lr_tag(39 downto 20),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(15 downto 8),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 2),
      memory_space_1_sr_req => memory_space_1_sr_req(1 downto 1),
      memory_space_1_sr_ack => memory_space_1_sr_ack(1 downto 1),
      memory_space_1_sr_addr => memory_space_1_sr_addr(1 downto 1),
      memory_space_1_sr_data => memory_space_1_sr_data(15 downto 8),
      memory_space_1_sr_tag => memory_space_1_sr_tag(39 downto 20),
      memory_space_1_sc_req => memory_space_1_sc_req(1 downto 1),
      memory_space_1_sc_ack => memory_space_1_sc_ack(1 downto 1),
      memory_space_1_sc_tag => memory_space_1_sc_tag(3 downto 2),
      tag_in => bz_tag_in,
      tag_out => bz_tag_out-- 
    ); -- 
  -- module call
  call_rs1_data <= call_in_args(79 downto 48);
  call_rs2_data <= call_in_args(47 downto 16);
  call_rd <= call_in_args(15 downto 8);
  call_pc <= call_in_args(7 downto 0);
  call_out_args <= call_next_pc ;
  -- call arbiter for module call
  call_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 80,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => call_call_reqs,
      call_acks => call_call_acks,
      return_reqs => call_return_reqs,
      return_acks => call_return_acks,
      call_data  => call_call_data,
      call_tag  => call_call_tag,
      return_tag  => call_return_tag,
      call_mtag => call_tag_in,
      return_mtag => call_tag_out,
      return_data =>call_return_data,
      call_mreq => call_start_req,
      call_mack => call_start_ack,
      return_mreq => call_fin_req,
      return_mack => call_fin_ack,
      call_mdata => call_in_args,
      return_mdata => call_out_args,
      clk => clk, 
      reset => reset --
    ); --
  call_instance:call-- 
    generic map(tag_length => 2)
    port map(-- 
      rs1_data => call_rs1_data,
      rs2_data => call_rs2_data,
      rd => call_rd,
      pc => call_pc,
      next_pc => call_next_pc,
      start_req => call_start_req,
      start_ack => call_start_ack,
      fin_req => call_fin_req,
      fin_ack => call_fin_ack,
      clk => clk,
      reset => reset,
      accessreg_call_reqs => accessreg_call_reqs(8 downto 8),
      accessreg_call_acks => accessreg_call_acks(8 downto 8),
      accessreg_call_data => accessreg_call_data(368 downto 328),
      accessreg_call_tag => accessreg_call_tag(17 downto 16),
      accessreg_return_reqs => accessreg_return_reqs(8 downto 8),
      accessreg_return_acks => accessreg_return_acks(8 downto 8),
      accessreg_return_data => accessreg_return_data(287 downto 256),
      accessreg_return_tag => accessreg_return_tag(17 downto 16),
      tag_in => call_tag_in,
      tag_out => call_tag_out-- 
    ); -- 
  -- module cmp
  cmp_rs1_data <= cmp_in_args(79 downto 48);
  cmp_rs2_data <= cmp_in_args(47 downto 16);
  cmp_rd <= cmp_in_args(15 downto 8);
  cmp_pc <= cmp_in_args(7 downto 0);
  cmp_out_args <= cmp_next_pc ;
  -- call arbiter for module cmp
  cmp_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 80,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => cmp_call_reqs,
      call_acks => cmp_call_acks,
      return_reqs => cmp_return_reqs,
      return_acks => cmp_return_acks,
      call_data  => cmp_call_data,
      call_tag  => cmp_call_tag,
      return_tag  => cmp_return_tag,
      call_mtag => cmp_tag_in,
      return_mtag => cmp_tag_out,
      return_data =>cmp_return_data,
      call_mreq => cmp_start_req,
      call_mack => cmp_start_ack,
      return_mreq => cmp_fin_req,
      return_mack => cmp_fin_ack,
      call_mdata => cmp_in_args,
      return_mdata => cmp_out_args,
      clk => clk, 
      reset => reset --
    ); --
  cmp_instance:cmp-- 
    generic map(tag_length => 2)
    port map(-- 
      rs1_data => cmp_rs1_data,
      rs2_data => cmp_rs2_data,
      rd => cmp_rd,
      pc => cmp_pc,
      next_pc => cmp_next_pc,
      start_req => cmp_start_req,
      start_ack => cmp_start_ack,
      fin_req => cmp_fin_req,
      fin_ack => cmp_fin_ack,
      clk => clk,
      reset => reset,
      accessreg_call_reqs => accessreg_call_reqs(13 downto 13),
      accessreg_call_acks => accessreg_call_acks(13 downto 13),
      accessreg_call_data => accessreg_call_data(573 downto 533),
      accessreg_call_tag => accessreg_call_tag(27 downto 26),
      accessreg_return_reqs => accessreg_return_reqs(13 downto 13),
      accessreg_return_acks => accessreg_return_acks(13 downto 13),
      accessreg_return_data => accessreg_return_data(447 downto 416),
      accessreg_return_tag => accessreg_return_tag(27 downto 26),
      tag_in => cmp_tag_in,
      tag_out => cmp_tag_out-- 
    ); -- 
  -- module halt
  halt_pc <= halt_in_args(7 downto 0);
  halt_out_args <= halt_next_pc ;
  -- call arbiter for module halt
  halt_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 8,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => halt_call_reqs,
      call_acks => halt_call_acks,
      return_reqs => halt_return_reqs,
      return_acks => halt_return_acks,
      call_data  => halt_call_data,
      call_tag  => halt_call_tag,
      return_tag  => halt_return_tag,
      call_mtag => halt_tag_in,
      return_mtag => halt_tag_out,
      return_data =>halt_return_data,
      call_mreq => halt_start_req,
      call_mack => halt_start_ack,
      return_mreq => halt_fin_req,
      return_mack => halt_fin_ack,
      call_mdata => halt_in_args,
      return_mdata => halt_out_args,
      clk => clk, 
      reset => reset --
    ); --
  halt_instance:halt-- 
    generic map(tag_length => 2)
    port map(-- 
      pc => halt_pc,
      next_pc => halt_next_pc,
      start_req => halt_start_req,
      start_ack => halt_start_ack,
      fin_req => halt_fin_req,
      fin_ack => halt_fin_ack,
      clk => clk,
      reset => reset,
      tag_in => halt_tag_in,
      tag_out => halt_tag_out-- 
    ); -- 
  -- module init_mem
  -- call arbiter for module init_mem
  init_mem_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => init_mem_call_reqs,
      call_acks => init_mem_call_acks,
      return_reqs => init_mem_return_reqs,
      return_acks => init_mem_return_acks,
      call_tag  => init_mem_call_tag,
      return_tag  => init_mem_return_tag,
      call_mtag => init_mem_tag_in,
      return_mtag => init_mem_tag_out,
      call_mreq => init_mem_start_req,
      call_mack => init_mem_start_ack,
      return_mreq => init_mem_fin_req,
      return_mack => init_mem_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  init_mem_instance:init_mem-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => init_mem_start_req,
      start_ack => init_mem_start_ack,
      fin_req => init_mem_fin_req,
      fin_ack => init_mem_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(7 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(31 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(17 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(0 downto 0),
      tag_in => init_mem_tag_in,
      tag_out => init_mem_tag_out-- 
    ); -- 
  -- module init_reg
  -- call arbiter for module init_reg
  init_reg_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => init_reg_call_reqs,
      call_acks => init_reg_call_acks,
      return_reqs => init_reg_return_reqs,
      return_acks => init_reg_return_acks,
      call_tag  => init_reg_call_tag,
      return_tag  => init_reg_return_tag,
      call_mtag => init_reg_tag_in,
      return_mtag => init_reg_tag_out,
      call_mreq => init_reg_start_req,
      call_mack => init_reg_start_ack,
      return_mreq => init_reg_fin_req,
      return_mack => init_reg_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  init_reg_instance:init_reg-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => init_reg_start_req,
      start_ack => init_reg_start_ack,
      fin_req => init_reg_fin_req,
      fin_ack => init_reg_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(7 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(31 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(17 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      tag_in => init_reg_tag_in,
      tag_out => init_reg_tag_out-- 
    ); -- 
  -- module jmp
  jmp_rs1_data <= jmp_in_args(39 downto 8);
  jmp_pc <= jmp_in_args(7 downto 0);
  jmp_out_args <= jmp_next_pc ;
  -- call arbiter for module jmp
  jmp_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 40,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => jmp_call_reqs,
      call_acks => jmp_call_acks,
      return_reqs => jmp_return_reqs,
      return_acks => jmp_return_acks,
      call_data  => jmp_call_data,
      call_tag  => jmp_call_tag,
      return_tag  => jmp_return_tag,
      call_mtag => jmp_tag_in,
      return_mtag => jmp_tag_out,
      return_data =>jmp_return_data,
      call_mreq => jmp_start_req,
      call_mack => jmp_start_ack,
      return_mreq => jmp_fin_req,
      return_mack => jmp_fin_ack,
      call_mdata => jmp_in_args,
      return_mdata => jmp_out_args,
      clk => clk, 
      reset => reset --
    ); --
  jmp_instance:jmp-- 
    generic map(tag_length => 2)
    port map(-- 
      rs1_data => jmp_rs1_data,
      pc => jmp_pc,
      next_pc => jmp_next_pc,
      start_req => jmp_start_req,
      start_ack => jmp_start_ack,
      fin_req => jmp_fin_req,
      fin_ack => jmp_fin_ack,
      clk => clk,
      reset => reset,
      tag_in => jmp_tag_in,
      tag_out => jmp_tag_out-- 
    ); -- 
  -- module load
  load_rs1_data <= load_in_args(47 downto 16);
  load_rd <= load_in_args(15 downto 8);
  load_pc <= load_in_args(7 downto 0);
  load_out_args <= load_next_pc ;
  -- call arbiter for module load
  load_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 48,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => load_call_reqs,
      call_acks => load_call_acks,
      return_reqs => load_return_reqs,
      return_acks => load_return_acks,
      call_data  => load_call_data,
      call_tag  => load_call_tag,
      return_tag  => load_return_tag,
      call_mtag => load_tag_in,
      return_mtag => load_tag_out,
      return_data =>load_return_data,
      call_mreq => load_start_req,
      call_mack => load_start_ack,
      return_mreq => load_fin_req,
      return_mack => load_fin_ack,
      call_mdata => load_in_args,
      return_mdata => load_out_args,
      clk => clk, 
      reset => reset --
    ); --
  load_instance:load-- 
    generic map(tag_length => 2)
    port map(-- 
      rs1_data => load_rs1_data,
      rd => load_rd,
      pc => load_pc,
      next_pc => load_next_pc,
      start_req => load_start_req,
      start_ack => load_start_ack,
      fin_req => load_fin_req,
      fin_ack => load_fin_ack,
      clk => clk,
      reset => reset,
      accessMem_call_reqs => accessMem_call_reqs(1 downto 1),
      accessMem_call_acks => accessMem_call_acks(1 downto 1),
      accessMem_call_data => accessMem_call_data(81 downto 41),
      accessMem_call_tag => accessMem_call_tag(1 downto 1),
      accessMem_return_reqs => accessMem_return_reqs(1 downto 1),
      accessMem_return_acks => accessMem_return_acks(1 downto 1),
      accessMem_return_data => accessMem_return_data(63 downto 32),
      accessMem_return_tag => accessMem_return_tag(1 downto 1),
      accessreg_call_reqs => accessreg_call_reqs(3 downto 3),
      accessreg_call_acks => accessreg_call_acks(3 downto 3),
      accessreg_call_data => accessreg_call_data(163 downto 123),
      accessreg_call_tag => accessreg_call_tag(7 downto 6),
      accessreg_return_reqs => accessreg_return_reqs(3 downto 3),
      accessreg_return_acks => accessreg_return_acks(3 downto 3),
      accessreg_return_data => accessreg_return_data(127 downto 96),
      accessreg_return_tag => accessreg_return_tag(7 downto 6),
      tag_in => load_tag_in,
      tag_out => load_tag_out-- 
    ); -- 
  -- module or_i
  or_i_rs1_data <= or_i_in_args(79 downto 48);
  or_i_rs2_data <= or_i_in_args(47 downto 16);
  or_i_rd <= or_i_in_args(15 downto 8);
  or_i_pc <= or_i_in_args(7 downto 0);
  or_i_out_args <= or_i_next_pc ;
  -- call arbiter for module or_i
  or_i_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 80,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => or_i_call_reqs,
      call_acks => or_i_call_acks,
      return_reqs => or_i_return_reqs,
      return_acks => or_i_return_acks,
      call_data  => or_i_call_data,
      call_tag  => or_i_call_tag,
      return_tag  => or_i_return_tag,
      call_mtag => or_i_tag_in,
      return_mtag => or_i_tag_out,
      return_data =>or_i_return_data,
      call_mreq => or_i_start_req,
      call_mack => or_i_start_ack,
      return_mreq => or_i_fin_req,
      return_mack => or_i_fin_ack,
      call_mdata => or_i_in_args,
      return_mdata => or_i_out_args,
      clk => clk, 
      reset => reset --
    ); --
  or_i_instance:or_i-- 
    generic map(tag_length => 2)
    port map(-- 
      rs1_data => or_i_rs1_data,
      rs2_data => or_i_rs2_data,
      rd => or_i_rd,
      pc => or_i_pc,
      next_pc => or_i_next_pc,
      start_req => or_i_start_req,
      start_ack => or_i_start_ack,
      fin_req => or_i_fin_req,
      fin_ack => or_i_fin_ack,
      clk => clk,
      reset => reset,
      accessreg_call_reqs => accessreg_call_reqs(4 downto 4),
      accessreg_call_acks => accessreg_call_acks(4 downto 4),
      accessreg_call_data => accessreg_call_data(204 downto 164),
      accessreg_call_tag => accessreg_call_tag(9 downto 8),
      accessreg_return_reqs => accessreg_return_reqs(4 downto 4),
      accessreg_return_acks => accessreg_return_acks(4 downto 4),
      accessreg_return_data => accessreg_return_data(159 downto 128),
      accessreg_return_tag => accessreg_return_tag(9 downto 8),
      tag_in => or_i_tag_in,
      tag_out => or_i_tag_out-- 
    ); -- 
  -- module sbir
  sbir_imm <= sbir_in_args(23 downto 16);
  sbir_rd <= sbir_in_args(15 downto 8);
  sbir_pc <= sbir_in_args(7 downto 0);
  sbir_out_args <= sbir_next_pc ;
  -- call arbiter for module sbir
  sbir_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 24,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sbir_call_reqs,
      call_acks => sbir_call_acks,
      return_reqs => sbir_return_reqs,
      return_acks => sbir_return_acks,
      call_data  => sbir_call_data,
      call_tag  => sbir_call_tag,
      return_tag  => sbir_return_tag,
      call_mtag => sbir_tag_in,
      return_mtag => sbir_tag_out,
      return_data =>sbir_return_data,
      call_mreq => sbir_start_req,
      call_mack => sbir_start_ack,
      return_mreq => sbir_fin_req,
      return_mack => sbir_fin_ack,
      call_mdata => sbir_in_args,
      return_mdata => sbir_out_args,
      clk => clk, 
      reset => reset --
    ); --
  sbir_instance:sbir-- 
    generic map(tag_length => 2)
    port map(-- 
      imm => sbir_imm,
      rd => sbir_rd,
      pc => sbir_pc,
      next_pc => sbir_next_pc,
      start_req => sbir_start_req,
      start_ack => sbir_start_ack,
      fin_req => sbir_fin_req,
      fin_ack => sbir_fin_ack,
      clk => clk,
      reset => reset,
      accessreg_call_reqs => accessreg_call_reqs(5 downto 5),
      accessreg_call_acks => accessreg_call_acks(5 downto 5),
      accessreg_call_data => accessreg_call_data(245 downto 205),
      accessreg_call_tag => accessreg_call_tag(11 downto 10),
      accessreg_return_reqs => accessreg_return_reqs(5 downto 5),
      accessreg_return_acks => accessreg_return_acks(5 downto 5),
      accessreg_return_data => accessreg_return_data(191 downto 160),
      accessreg_return_tag => accessreg_return_tag(11 downto 10),
      tag_in => sbir_tag_in,
      tag_out => sbir_tag_out-- 
    ); -- 
  -- module sll_i
  sll_i_rs1_data <= sll_i_in_args(79 downto 48);
  sll_i_rs2_data <= sll_i_in_args(47 downto 16);
  sll_i_rd <= sll_i_in_args(15 downto 8);
  sll_i_pc <= sll_i_in_args(7 downto 0);
  sll_i_out_args <= sll_i_next_pc ;
  -- call arbiter for module sll_i
  sll_i_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 80,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sll_i_call_reqs,
      call_acks => sll_i_call_acks,
      return_reqs => sll_i_return_reqs,
      return_acks => sll_i_return_acks,
      call_data  => sll_i_call_data,
      call_tag  => sll_i_call_tag,
      return_tag  => sll_i_return_tag,
      call_mtag => sll_i_tag_in,
      return_mtag => sll_i_tag_out,
      return_data =>sll_i_return_data,
      call_mreq => sll_i_start_req,
      call_mack => sll_i_start_ack,
      return_mreq => sll_i_fin_req,
      return_mack => sll_i_fin_ack,
      call_mdata => sll_i_in_args,
      return_mdata => sll_i_out_args,
      clk => clk, 
      reset => reset --
    ); --
  sll_i_instance:sll_i-- 
    generic map(tag_length => 2)
    port map(-- 
      rs1_data => sll_i_rs1_data,
      rs2_data => sll_i_rs2_data,
      rd => sll_i_rd,
      pc => sll_i_pc,
      next_pc => sll_i_next_pc,
      start_req => sll_i_start_req,
      start_ack => sll_i_start_ack,
      fin_req => sll_i_fin_req,
      fin_ack => sll_i_fin_ack,
      clk => clk,
      reset => reset,
      accessreg_call_reqs => accessreg_call_reqs(10 downto 10),
      accessreg_call_acks => accessreg_call_acks(10 downto 10),
      accessreg_call_data => accessreg_call_data(450 downto 410),
      accessreg_call_tag => accessreg_call_tag(21 downto 20),
      accessreg_return_reqs => accessreg_return_reqs(10 downto 10),
      accessreg_return_acks => accessreg_return_acks(10 downto 10),
      accessreg_return_data => accessreg_return_data(351 downto 320),
      accessreg_return_tag => accessreg_return_tag(21 downto 20),
      tag_in => sll_i_tag_in,
      tag_out => sll_i_tag_out-- 
    ); -- 
  -- module sra_i
  sra_i_rs1_data <= sra_i_in_args(79 downto 48);
  sra_i_rs2_data <= sra_i_in_args(47 downto 16);
  sra_i_rd <= sra_i_in_args(15 downto 8);
  sra_i_pc <= sra_i_in_args(7 downto 0);
  sra_i_out_args <= sra_i_next_pc ;
  -- call arbiter for module sra_i
  sra_i_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 80,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sra_i_call_reqs,
      call_acks => sra_i_call_acks,
      return_reqs => sra_i_return_reqs,
      return_acks => sra_i_return_acks,
      call_data  => sra_i_call_data,
      call_tag  => sra_i_call_tag,
      return_tag  => sra_i_return_tag,
      call_mtag => sra_i_tag_in,
      return_mtag => sra_i_tag_out,
      return_data =>sra_i_return_data,
      call_mreq => sra_i_start_req,
      call_mack => sra_i_start_ack,
      return_mreq => sra_i_fin_req,
      return_mack => sra_i_fin_ack,
      call_mdata => sra_i_in_args,
      return_mdata => sra_i_out_args,
      clk => clk, 
      reset => reset --
    ); --
  sra_i_instance:sra_i-- 
    generic map(tag_length => 2)
    port map(-- 
      rs1_data => sra_i_rs1_data,
      rs2_data => sra_i_rs2_data,
      rd => sra_i_rd,
      pc => sra_i_pc,
      next_pc => sra_i_next_pc,
      start_req => sra_i_start_req,
      start_ack => sra_i_start_ack,
      fin_req => sra_i_fin_req,
      fin_ack => sra_i_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(0 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(19 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(31 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(2 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(0 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(31 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(19 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(2 downto 0),
      accessreg_call_reqs => accessreg_call_reqs(6 downto 6),
      accessreg_call_acks => accessreg_call_acks(6 downto 6),
      accessreg_call_data => accessreg_call_data(286 downto 246),
      accessreg_call_tag => accessreg_call_tag(13 downto 12),
      accessreg_return_reqs => accessreg_return_reqs(6 downto 6),
      accessreg_return_acks => accessreg_return_acks(6 downto 6),
      accessreg_return_data => accessreg_return_data(223 downto 192),
      accessreg_return_tag => accessreg_return_tag(13 downto 12),
      tag_in => sra_i_tag_in,
      tag_out => sra_i_tag_out-- 
    ); -- 
  -- module srl_i
  srl_i_rs1_data <= srl_i_in_args(79 downto 48);
  srl_i_rs2_data <= srl_i_in_args(47 downto 16);
  srl_i_rd <= srl_i_in_args(15 downto 8);
  srl_i_pc <= srl_i_in_args(7 downto 0);
  srl_i_out_args <= srl_i_next_pc ;
  -- call arbiter for module srl_i
  srl_i_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 80,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => srl_i_call_reqs,
      call_acks => srl_i_call_acks,
      return_reqs => srl_i_return_reqs,
      return_acks => srl_i_return_acks,
      call_data  => srl_i_call_data,
      call_tag  => srl_i_call_tag,
      return_tag  => srl_i_return_tag,
      call_mtag => srl_i_tag_in,
      return_mtag => srl_i_tag_out,
      return_data =>srl_i_return_data,
      call_mreq => srl_i_start_req,
      call_mack => srl_i_start_ack,
      return_mreq => srl_i_fin_req,
      return_mack => srl_i_fin_ack,
      call_mdata => srl_i_in_args,
      return_mdata => srl_i_out_args,
      clk => clk, 
      reset => reset --
    ); --
  srl_i_instance:srl_i-- 
    generic map(tag_length => 2)
    port map(-- 
      rs1_data => srl_i_rs1_data,
      rs2_data => srl_i_rs2_data,
      rd => srl_i_rd,
      pc => srl_i_pc,
      next_pc => srl_i_next_pc,
      start_req => srl_i_start_req,
      start_ack => srl_i_start_ack,
      fin_req => srl_i_fin_req,
      fin_ack => srl_i_fin_ack,
      clk => clk,
      reset => reset,
      accessreg_call_reqs => accessreg_call_reqs(2 downto 2),
      accessreg_call_acks => accessreg_call_acks(2 downto 2),
      accessreg_call_data => accessreg_call_data(122 downto 82),
      accessreg_call_tag => accessreg_call_tag(5 downto 4),
      accessreg_return_reqs => accessreg_return_reqs(2 downto 2),
      accessreg_return_acks => accessreg_return_acks(2 downto 2),
      accessreg_return_data => accessreg_return_data(95 downto 64),
      accessreg_return_tag => accessreg_return_tag(5 downto 4),
      tag_in => srl_i_tag_in,
      tag_out => srl_i_tag_out-- 
    ); -- 
  -- module store
  store_rs1_data <= store_in_args(71 downto 40);
  store_rs2_data <= store_in_args(39 downto 8);
  store_pc <= store_in_args(7 downto 0);
  store_out_args <= store_next_pc ;
  -- call arbiter for module store
  store_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 72,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => store_call_reqs,
      call_acks => store_call_acks,
      return_reqs => store_return_reqs,
      return_acks => store_return_acks,
      call_data  => store_call_data,
      call_tag  => store_call_tag,
      return_tag  => store_return_tag,
      call_mtag => store_tag_in,
      return_mtag => store_tag_out,
      return_data =>store_return_data,
      call_mreq => store_start_req,
      call_mack => store_start_ack,
      return_mreq => store_fin_req,
      return_mack => store_fin_ack,
      call_mdata => store_in_args,
      return_mdata => store_out_args,
      clk => clk, 
      reset => reset --
    ); --
  store_instance:store-- 
    generic map(tag_length => 2)
    port map(-- 
      rs1_data => store_rs1_data,
      rs2_data => store_rs2_data,
      pc => store_pc,
      next_pc => store_next_pc,
      start_req => store_start_req,
      start_ack => store_start_ack,
      fin_req => store_fin_req,
      fin_ack => store_fin_ack,
      clk => clk,
      reset => reset,
      accessMem_call_reqs => accessMem_call_reqs(0 downto 0),
      accessMem_call_acks => accessMem_call_acks(0 downto 0),
      accessMem_call_data => accessMem_call_data(40 downto 0),
      accessMem_call_tag => accessMem_call_tag(0 downto 0),
      accessMem_return_reqs => accessMem_return_reqs(0 downto 0),
      accessMem_return_acks => accessMem_return_acks(0 downto 0),
      accessMem_return_data => accessMem_return_data(31 downto 0),
      accessMem_return_tag => accessMem_return_tag(0 downto 0),
      tag_in => store_tag_in,
      tag_out => store_tag_out-- 
    ); -- 
  -- module sub
  sub_rs1_data <= sub_in_args(79 downto 48);
  sub_rs2_data <= sub_in_args(47 downto 16);
  sub_rd <= sub_in_args(15 downto 8);
  sub_pc <= sub_in_args(7 downto 0);
  sub_out_args <= sub_next_pc ;
  -- call arbiter for module sub
  sub_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 80,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sub_call_reqs,
      call_acks => sub_call_acks,
      return_reqs => sub_return_reqs,
      return_acks => sub_return_acks,
      call_data  => sub_call_data,
      call_tag  => sub_call_tag,
      return_tag  => sub_return_tag,
      call_mtag => sub_tag_in,
      return_mtag => sub_tag_out,
      return_data =>sub_return_data,
      call_mreq => sub_start_req,
      call_mack => sub_start_ack,
      return_mreq => sub_fin_req,
      return_mack => sub_fin_ack,
      call_mdata => sub_in_args,
      return_mdata => sub_out_args,
      clk => clk, 
      reset => reset --
    ); --
  sub_instance:sub-- 
    generic map(tag_length => 2)
    port map(-- 
      rs1_data => sub_rs1_data,
      rs2_data => sub_rs2_data,
      rd => sub_rd,
      pc => sub_pc,
      next_pc => sub_next_pc,
      start_req => sub_start_req,
      start_ack => sub_start_ack,
      fin_req => sub_fin_req,
      fin_ack => sub_fin_ack,
      clk => clk,
      reset => reset,
      accessreg_call_reqs => accessreg_call_reqs(12 downto 12),
      accessreg_call_acks => accessreg_call_acks(12 downto 12),
      accessreg_call_data => accessreg_call_data(532 downto 492),
      accessreg_call_tag => accessreg_call_tag(25 downto 24),
      accessreg_return_reqs => accessreg_return_reqs(12 downto 12),
      accessreg_return_acks => accessreg_return_acks(12 downto 12),
      accessreg_return_data => accessreg_return_data(415 downto 384),
      accessreg_return_tag => accessreg_return_tag(25 downto 24),
      tag_in => sub_tag_in,
      tag_out => sub_tag_out-- 
    ); -- 
  -- module try
  try_pc <= try_in_args(39 downto 32);
  try_inst <= try_in_args(31 downto 0);
  try_out_args <= try_next_pc ;
  -- call arbiter for module try
  try_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 40,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => try_call_reqs,
      call_acks => try_call_acks,
      return_reqs => try_return_reqs,
      return_acks => try_return_acks,
      call_data  => try_call_data,
      call_tag  => try_call_tag,
      return_tag  => try_return_tag,
      call_mtag => try_tag_in,
      return_mtag => try_tag_out,
      return_data =>try_return_data,
      call_mreq => try_start_req,
      call_mack => try_start_ack,
      return_mreq => try_fin_req,
      return_mack => try_fin_ack,
      call_mdata => try_in_args,
      return_mdata => try_out_args,
      clk => clk, 
      reset => reset --
    ); --
  try_instance:try-- 
    generic map(tag_length => 2)
    port map(-- 
      pc => try_pc,
      inst => try_inst,
      next_pc => try_next_pc,
      start_req => try_start_req,
      start_ack => try_start_ack,
      fin_req => try_fin_req,
      fin_ack => try_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(0 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(19 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(7 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(0 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(7 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(19 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(1 downto 0),
      accessreg_call_reqs => accessreg_call_reqs(0 downto 0),
      accessreg_call_acks => accessreg_call_acks(0 downto 0),
      accessreg_call_data => accessreg_call_data(40 downto 0),
      accessreg_call_tag => accessreg_call_tag(1 downto 0),
      accessreg_return_reqs => accessreg_return_reqs(0 downto 0),
      accessreg_return_acks => accessreg_return_acks(0 downto 0),
      accessreg_return_data => accessreg_return_data(31 downto 0),
      accessreg_return_tag => accessreg_return_tag(1 downto 0),
      add_call_reqs => add_call_reqs(0 downto 0),
      add_call_acks => add_call_acks(0 downto 0),
      add_call_data => add_call_data(79 downto 0),
      add_call_tag => add_call_tag(0 downto 0),
      add_return_reqs => add_return_reqs(0 downto 0),
      add_return_acks => add_return_acks(0 downto 0),
      add_return_data => add_return_data(7 downto 0),
      add_return_tag => add_return_tag(0 downto 0),
      and_i_call_reqs => and_i_call_reqs(0 downto 0),
      and_i_call_acks => and_i_call_acks(0 downto 0),
      and_i_call_data => and_i_call_data(79 downto 0),
      and_i_call_tag => and_i_call_tag(0 downto 0),
      and_i_return_reqs => and_i_return_reqs(0 downto 0),
      and_i_return_acks => and_i_return_acks(0 downto 0),
      and_i_return_data => and_i_return_data(7 downto 0),
      and_i_return_tag => and_i_return_tag(0 downto 0),
      bn_call_reqs => bn_call_reqs(0 downto 0),
      bn_call_acks => bn_call_acks(0 downto 0),
      bn_call_data => bn_call_data(79 downto 0),
      bn_call_tag => bn_call_tag(0 downto 0),
      bn_return_reqs => bn_return_reqs(0 downto 0),
      bn_return_acks => bn_return_acks(0 downto 0),
      bn_return_data => bn_return_data(7 downto 0),
      bn_return_tag => bn_return_tag(0 downto 0),
      bz_call_reqs => bz_call_reqs(0 downto 0),
      bz_call_acks => bz_call_acks(0 downto 0),
      bz_call_data => bz_call_data(79 downto 0),
      bz_call_tag => bz_call_tag(0 downto 0),
      bz_return_reqs => bz_return_reqs(0 downto 0),
      bz_return_acks => bz_return_acks(0 downto 0),
      bz_return_data => bz_return_data(7 downto 0),
      bz_return_tag => bz_return_tag(0 downto 0),
      call_call_reqs => call_call_reqs(0 downto 0),
      call_call_acks => call_call_acks(0 downto 0),
      call_call_data => call_call_data(79 downto 0),
      call_call_tag => call_call_tag(0 downto 0),
      call_return_reqs => call_return_reqs(0 downto 0),
      call_return_acks => call_return_acks(0 downto 0),
      call_return_data => call_return_data(7 downto 0),
      call_return_tag => call_return_tag(0 downto 0),
      cmp_call_reqs => cmp_call_reqs(0 downto 0),
      cmp_call_acks => cmp_call_acks(0 downto 0),
      cmp_call_data => cmp_call_data(79 downto 0),
      cmp_call_tag => cmp_call_tag(0 downto 0),
      cmp_return_reqs => cmp_return_reqs(0 downto 0),
      cmp_return_acks => cmp_return_acks(0 downto 0),
      cmp_return_data => cmp_return_data(7 downto 0),
      cmp_return_tag => cmp_return_tag(0 downto 0),
      halt_call_reqs => halt_call_reqs(0 downto 0),
      halt_call_acks => halt_call_acks(0 downto 0),
      halt_call_data => halt_call_data(7 downto 0),
      halt_call_tag => halt_call_tag(0 downto 0),
      halt_return_reqs => halt_return_reqs(0 downto 0),
      halt_return_acks => halt_return_acks(0 downto 0),
      halt_return_data => halt_return_data(7 downto 0),
      halt_return_tag => halt_return_tag(0 downto 0),
      jmp_call_reqs => jmp_call_reqs(0 downto 0),
      jmp_call_acks => jmp_call_acks(0 downto 0),
      jmp_call_data => jmp_call_data(39 downto 0),
      jmp_call_tag => jmp_call_tag(0 downto 0),
      jmp_return_reqs => jmp_return_reqs(0 downto 0),
      jmp_return_acks => jmp_return_acks(0 downto 0),
      jmp_return_data => jmp_return_data(7 downto 0),
      jmp_return_tag => jmp_return_tag(0 downto 0),
      load_call_reqs => load_call_reqs(0 downto 0),
      load_call_acks => load_call_acks(0 downto 0),
      load_call_data => load_call_data(47 downto 0),
      load_call_tag => load_call_tag(0 downto 0),
      load_return_reqs => load_return_reqs(0 downto 0),
      load_return_acks => load_return_acks(0 downto 0),
      load_return_data => load_return_data(7 downto 0),
      load_return_tag => load_return_tag(0 downto 0),
      or_i_call_reqs => or_i_call_reqs(0 downto 0),
      or_i_call_acks => or_i_call_acks(0 downto 0),
      or_i_call_data => or_i_call_data(79 downto 0),
      or_i_call_tag => or_i_call_tag(0 downto 0),
      or_i_return_reqs => or_i_return_reqs(0 downto 0),
      or_i_return_acks => or_i_return_acks(0 downto 0),
      or_i_return_data => or_i_return_data(7 downto 0),
      or_i_return_tag => or_i_return_tag(0 downto 0),
      sbir_call_reqs => sbir_call_reqs(0 downto 0),
      sbir_call_acks => sbir_call_acks(0 downto 0),
      sbir_call_data => sbir_call_data(23 downto 0),
      sbir_call_tag => sbir_call_tag(0 downto 0),
      sbir_return_reqs => sbir_return_reqs(0 downto 0),
      sbir_return_acks => sbir_return_acks(0 downto 0),
      sbir_return_data => sbir_return_data(7 downto 0),
      sbir_return_tag => sbir_return_tag(0 downto 0),
      sll_i_call_reqs => sll_i_call_reqs(0 downto 0),
      sll_i_call_acks => sll_i_call_acks(0 downto 0),
      sll_i_call_data => sll_i_call_data(79 downto 0),
      sll_i_call_tag => sll_i_call_tag(0 downto 0),
      sll_i_return_reqs => sll_i_return_reqs(0 downto 0),
      sll_i_return_acks => sll_i_return_acks(0 downto 0),
      sll_i_return_data => sll_i_return_data(7 downto 0),
      sll_i_return_tag => sll_i_return_tag(0 downto 0),
      sra_i_call_reqs => sra_i_call_reqs(0 downto 0),
      sra_i_call_acks => sra_i_call_acks(0 downto 0),
      sra_i_call_data => sra_i_call_data(79 downto 0),
      sra_i_call_tag => sra_i_call_tag(0 downto 0),
      sra_i_return_reqs => sra_i_return_reqs(0 downto 0),
      sra_i_return_acks => sra_i_return_acks(0 downto 0),
      sra_i_return_data => sra_i_return_data(7 downto 0),
      sra_i_return_tag => sra_i_return_tag(0 downto 0),
      srl_i_call_reqs => srl_i_call_reqs(0 downto 0),
      srl_i_call_acks => srl_i_call_acks(0 downto 0),
      srl_i_call_data => srl_i_call_data(79 downto 0),
      srl_i_call_tag => srl_i_call_tag(0 downto 0),
      srl_i_return_reqs => srl_i_return_reqs(0 downto 0),
      srl_i_return_acks => srl_i_return_acks(0 downto 0),
      srl_i_return_data => srl_i_return_data(7 downto 0),
      srl_i_return_tag => srl_i_return_tag(0 downto 0),
      store_call_reqs => store_call_reqs(0 downto 0),
      store_call_acks => store_call_acks(0 downto 0),
      store_call_data => store_call_data(71 downto 0),
      store_call_tag => store_call_tag(0 downto 0),
      store_return_reqs => store_return_reqs(0 downto 0),
      store_return_acks => store_return_acks(0 downto 0),
      store_return_data => store_return_data(7 downto 0),
      store_return_tag => store_return_tag(0 downto 0),
      sub_call_reqs => sub_call_reqs(0 downto 0),
      sub_call_acks => sub_call_acks(0 downto 0),
      sub_call_data => sub_call_data(79 downto 0),
      sub_call_tag => sub_call_tag(0 downto 0),
      sub_return_reqs => sub_return_reqs(0 downto 0),
      sub_return_acks => sub_return_acks(0 downto 0),
      sub_return_data => sub_return_data(7 downto 0),
      sub_return_tag => sub_return_tag(0 downto 0),
      xnor_i_call_reqs => xnor_i_call_reqs(0 downto 0),
      xnor_i_call_acks => xnor_i_call_acks(0 downto 0),
      xnor_i_call_data => xnor_i_call_data(79 downto 0),
      xnor_i_call_tag => xnor_i_call_tag(0 downto 0),
      xnor_i_return_reqs => xnor_i_return_reqs(0 downto 0),
      xnor_i_return_acks => xnor_i_return_acks(0 downto 0),
      xnor_i_return_data => xnor_i_return_data(7 downto 0),
      xnor_i_return_tag => xnor_i_return_tag(0 downto 0),
      xor_i_call_reqs => xor_i_call_reqs(0 downto 0),
      xor_i_call_acks => xor_i_call_acks(0 downto 0),
      xor_i_call_data => xor_i_call_data(79 downto 0),
      xor_i_call_tag => xor_i_call_tag(0 downto 0),
      xor_i_return_reqs => xor_i_return_reqs(0 downto 0),
      xor_i_return_acks => xor_i_return_acks(0 downto 0),
      xor_i_return_data => xor_i_return_data(7 downto 0),
      xor_i_return_tag => xor_i_return_tag(0 downto 0),
      tag_in => try_tag_in,
      tag_out => try_tag_out-- 
    ); -- 
  -- module try1
  try1_instance:try1-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => try1_start_req,
      start_ack => try1_start_ack,
      fin_req => try1_fin_req,
      fin_ack => try1_fin_ack,
      clk => clk,
      reset => reset,
      write_mem_pipe_read_req => write_mem_pipe_read_req(0 downto 0),
      write_mem_pipe_read_ack => write_mem_pipe_read_ack(0 downto 0),
      write_mem_pipe_read_data => write_mem_pipe_read_data(7 downto 0),
      LEDS_pipe_write_req => LEDS_pipe_write_req(0 downto 0),
      LEDS_pipe_write_ack => LEDS_pipe_write_ack(0 downto 0),
      LEDS_pipe_write_data => LEDS_pipe_write_data(15 downto 0),
      reg_output_pipe_write_req => reg_output_pipe_write_req(0 downto 0),
      reg_output_pipe_write_ack => reg_output_pipe_write_ack(0 downto 0),
      reg_output_pipe_write_data => reg_output_pipe_write_data(7 downto 0),
      init_mem_call_reqs => init_mem_call_reqs(0 downto 0),
      init_mem_call_acks => init_mem_call_acks(0 downto 0),
      init_mem_call_tag => init_mem_call_tag(0 downto 0),
      init_mem_return_reqs => init_mem_return_reqs(0 downto 0),
      init_mem_return_acks => init_mem_return_acks(0 downto 0),
      init_mem_return_tag => init_mem_return_tag(0 downto 0),
      init_reg_call_reqs => init_reg_call_reqs(0 downto 0),
      init_reg_call_acks => init_reg_call_acks(0 downto 0),
      init_reg_call_tag => init_reg_call_tag(0 downto 0),
      init_reg_return_reqs => init_reg_return_reqs(0 downto 0),
      init_reg_return_acks => init_reg_return_acks(0 downto 0),
      init_reg_return_tag => init_reg_return_tag(0 downto 0),
      try_call_reqs => try_call_reqs(0 downto 0),
      try_call_acks => try_call_acks(0 downto 0),
      try_call_data => try_call_data(39 downto 0),
      try_call_tag => try_call_tag(0 downto 0),
      try_return_reqs => try_return_reqs(0 downto 0),
      try_return_acks => try_return_acks(0 downto 0),
      try_return_data => try_return_data(7 downto 0),
      try_return_tag => try_return_tag(0 downto 0),
      tag_in => try1_tag_in,
      tag_out => try1_tag_out-- 
    ); -- 
  -- module will be run forever 
  try1_tag_in <= (others => '0');
  try1_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => try1_start_req, start_ack => try1_start_ack,  fin_req => try1_fin_req,  fin_ack => try1_fin_ack);
  -- module xnor_i
  xnor_i_rs1_data <= xnor_i_in_args(79 downto 48);
  xnor_i_rs2_data <= xnor_i_in_args(47 downto 16);
  xnor_i_rd <= xnor_i_in_args(15 downto 8);
  xnor_i_pc <= xnor_i_in_args(7 downto 0);
  xnor_i_out_args <= xnor_i_next_pc ;
  -- call arbiter for module xnor_i
  xnor_i_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 80,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => xnor_i_call_reqs,
      call_acks => xnor_i_call_acks,
      return_reqs => xnor_i_return_reqs,
      return_acks => xnor_i_return_acks,
      call_data  => xnor_i_call_data,
      call_tag  => xnor_i_call_tag,
      return_tag  => xnor_i_return_tag,
      call_mtag => xnor_i_tag_in,
      return_mtag => xnor_i_tag_out,
      return_data =>xnor_i_return_data,
      call_mreq => xnor_i_start_req,
      call_mack => xnor_i_start_ack,
      return_mreq => xnor_i_fin_req,
      return_mack => xnor_i_fin_ack,
      call_mdata => xnor_i_in_args,
      return_mdata => xnor_i_out_args,
      clk => clk, 
      reset => reset --
    ); --
  xnor_i_instance:xnor_i-- 
    generic map(tag_length => 2)
    port map(-- 
      rs1_data => xnor_i_rs1_data,
      rs2_data => xnor_i_rs2_data,
      rd => xnor_i_rd,
      pc => xnor_i_pc,
      next_pc => xnor_i_next_pc,
      start_req => xnor_i_start_req,
      start_ack => xnor_i_start_ack,
      fin_req => xnor_i_fin_req,
      fin_ack => xnor_i_fin_ack,
      clk => clk,
      reset => reset,
      accessreg_call_reqs => accessreg_call_reqs(7 downto 7),
      accessreg_call_acks => accessreg_call_acks(7 downto 7),
      accessreg_call_data => accessreg_call_data(327 downto 287),
      accessreg_call_tag => accessreg_call_tag(15 downto 14),
      accessreg_return_reqs => accessreg_return_reqs(7 downto 7),
      accessreg_return_acks => accessreg_return_acks(7 downto 7),
      accessreg_return_data => accessreg_return_data(255 downto 224),
      accessreg_return_tag => accessreg_return_tag(15 downto 14),
      tag_in => xnor_i_tag_in,
      tag_out => xnor_i_tag_out-- 
    ); -- 
  -- module xor_i
  xor_i_rs1_data <= xor_i_in_args(79 downto 48);
  xor_i_rs2_data <= xor_i_in_args(47 downto 16);
  xor_i_rd <= xor_i_in_args(15 downto 8);
  xor_i_pc <= xor_i_in_args(7 downto 0);
  xor_i_out_args <= xor_i_next_pc ;
  -- call arbiter for module xor_i
  xor_i_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 80,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => xor_i_call_reqs,
      call_acks => xor_i_call_acks,
      return_reqs => xor_i_return_reqs,
      return_acks => xor_i_return_acks,
      call_data  => xor_i_call_data,
      call_tag  => xor_i_call_tag,
      return_tag  => xor_i_return_tag,
      call_mtag => xor_i_tag_in,
      return_mtag => xor_i_tag_out,
      return_data =>xor_i_return_data,
      call_mreq => xor_i_start_req,
      call_mack => xor_i_start_ack,
      return_mreq => xor_i_fin_req,
      return_mack => xor_i_fin_ack,
      call_mdata => xor_i_in_args,
      return_mdata => xor_i_out_args,
      clk => clk, 
      reset => reset --
    ); --
  xor_i_instance:xor_i-- 
    generic map(tag_length => 2)
    port map(-- 
      rs1_data => xor_i_rs1_data,
      rs2_data => xor_i_rs2_data,
      rd => xor_i_rd,
      pc => xor_i_pc,
      next_pc => xor_i_next_pc,
      start_req => xor_i_start_req,
      start_ack => xor_i_start_ack,
      fin_req => xor_i_fin_req,
      fin_ack => xor_i_fin_ack,
      clk => clk,
      reset => reset,
      accessreg_call_reqs => accessreg_call_reqs(1 downto 1),
      accessreg_call_acks => accessreg_call_acks(1 downto 1),
      accessreg_call_data => accessreg_call_data(81 downto 41),
      accessreg_call_tag => accessreg_call_tag(3 downto 2),
      accessreg_return_reqs => accessreg_return_reqs(1 downto 1),
      accessreg_return_acks => accessreg_return_acks(1 downto 1),
      accessreg_return_data => accessreg_return_data(63 downto 32),
      accessreg_return_tag => accessreg_return_tag(3 downto 2),
      tag_in => xor_i_tag_in,
      tag_out => xor_i_tag_out-- 
    ); -- 
  LEDS_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe LEDS",
      volatile_flag => false,
      num_writes => 1,
      data_width => 16 --
    ) 
    port map( -- 
      read_data => LEDS,
      write_req => LEDS_pipe_write_req,
      write_ack => LEDS_pipe_write_ack,
      write_data => LEDS_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  reg_output_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe reg_output",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 40 --
    )
    port map( -- 
      read_req => reg_output_pipe_read_req,
      read_ack => reg_output_pipe_read_ack,
      read_data => reg_output_pipe_read_data,
      write_req => reg_output_pipe_write_req,
      write_ack => reg_output_pipe_write_ack,
      write_data => reg_output_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  write_mem_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe write_mem",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 40 --
    )
    port map( -- 
      read_req => write_mem_pipe_read_req,
      read_ack => write_mem_pipe_read_ack,
      read_data => write_mem_pipe_read_data,
      write_req => write_mem_pipe_write_req,
      write_ack => write_mem_pipe_write_ack,
      write_data => write_mem_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 2,
      addr_width => 8,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 8,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 3,
      num_stores => 3,
      addr_width => 1,
      data_width => 8,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 2,
      addr_width => 8,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 8,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
